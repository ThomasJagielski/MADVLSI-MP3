magic
tech sky130A
timestamp 1615609162
<< nmos >>
rect -15 -1765 35 -1165
rect 85 -1765 135 -1165
rect 185 -1765 235 -1165
rect 285 -1765 335 -1165
rect 385 -1765 435 -1165
rect 485 -1765 535 -1165
rect 585 -1765 635 -1165
rect 685 -1765 735 -1165
rect 785 -1765 835 -1165
rect 885 -1765 935 -1165
<< ndiff >>
rect -65 -1180 -15 -1165
rect -65 -1750 -50 -1180
rect -30 -1750 -15 -1180
rect -65 -1765 -15 -1750
rect 35 -1180 85 -1165
rect 35 -1750 50 -1180
rect 70 -1750 85 -1180
rect 35 -1765 85 -1750
rect 135 -1180 185 -1165
rect 135 -1750 150 -1180
rect 170 -1750 185 -1180
rect 135 -1765 185 -1750
rect 235 -1180 285 -1165
rect 235 -1750 250 -1180
rect 270 -1750 285 -1180
rect 235 -1765 285 -1750
rect 335 -1180 385 -1165
rect 335 -1750 350 -1180
rect 370 -1750 385 -1180
rect 335 -1765 385 -1750
rect 435 -1180 485 -1165
rect 435 -1750 450 -1180
rect 470 -1750 485 -1180
rect 435 -1765 485 -1750
rect 535 -1180 585 -1165
rect 535 -1750 550 -1180
rect 570 -1750 585 -1180
rect 535 -1765 585 -1750
rect 635 -1180 685 -1165
rect 635 -1750 650 -1180
rect 670 -1750 685 -1180
rect 635 -1765 685 -1750
rect 735 -1180 785 -1165
rect 735 -1750 750 -1180
rect 770 -1750 785 -1180
rect 735 -1765 785 -1750
rect 835 -1180 885 -1165
rect 835 -1750 850 -1180
rect 870 -1750 885 -1180
rect 835 -1765 885 -1750
rect 935 -1180 985 -1165
rect 935 -1750 950 -1180
rect 970 -1750 985 -1180
rect 935 -1765 985 -1750
<< ndiffc >>
rect -50 -1750 -30 -1180
rect 50 -1750 70 -1180
rect 150 -1750 170 -1180
rect 250 -1750 270 -1180
rect 350 -1750 370 -1180
rect 450 -1750 470 -1180
rect 550 -1750 570 -1180
rect 650 -1750 670 -1180
rect 750 -1750 770 -1180
rect 850 -1750 870 -1180
rect 950 -1750 970 -1180
<< psubdiff >>
rect -115 -1180 -65 -1165
rect -115 -1750 -100 -1180
rect -80 -1750 -65 -1180
rect -115 -1765 -65 -1750
rect 985 -1180 1035 -1165
rect 985 -1750 1000 -1180
rect 1020 -1750 1035 -1180
rect 985 -1765 1035 -1750
<< psubdiffcont >>
rect -100 -1750 -80 -1180
rect 1000 -1750 1020 -1180
<< poly >>
rect 450 -950 470 -935
rect 380 -960 540 -950
rect 380 -980 390 -960
rect 410 -965 510 -960
rect 410 -980 420 -965
rect 380 -990 420 -980
rect 500 -980 510 -965
rect 530 -980 540 -960
rect 500 -990 540 -980
rect -60 -1060 -20 -1050
rect -60 -1080 -50 -1060
rect -30 -1075 -20 -1060
rect -30 -1080 100 -1075
rect -60 -1090 100 -1080
rect 85 -1110 100 -1090
rect -60 -1125 -20 -1115
rect -60 -1145 -50 -1125
rect -30 -1140 -20 -1125
rect 85 -1125 835 -1110
rect -30 -1145 35 -1140
rect -60 -1155 35 -1145
rect -15 -1165 35 -1155
rect 85 -1165 135 -1125
rect 185 -1165 235 -1150
rect 285 -1165 335 -1150
rect 385 -1165 435 -1125
rect 485 -1165 535 -1125
rect 585 -1165 635 -1150
rect 685 -1165 735 -1150
rect 785 -1165 835 -1125
rect 940 -1125 980 -1115
rect 940 -1140 950 -1125
rect 885 -1145 950 -1140
rect 970 -1145 980 -1125
rect 885 -1155 980 -1145
rect 885 -1165 935 -1155
rect -15 -1780 35 -1765
rect 85 -1780 135 -1765
rect 185 -1800 235 -1765
rect 285 -1800 335 -1765
rect 385 -1780 435 -1765
rect 485 -1780 535 -1765
rect -65 -1805 -25 -1800
rect 185 -1805 335 -1800
rect 585 -1805 635 -1765
rect 685 -1805 735 -1765
rect 785 -1780 835 -1765
rect 885 -1780 935 -1765
rect -65 -1810 735 -1805
rect -65 -1830 -55 -1810
rect -35 -1820 735 -1810
rect -35 -1830 -25 -1820
rect -65 -1840 -25 -1830
<< polycont >>
rect 390 -980 410 -960
rect 510 -980 530 -960
rect -50 -1080 -30 -1060
rect -50 -1145 -30 -1125
rect 950 -1145 970 -1125
rect -55 -1830 -35 -1810
<< locali >>
rect 40 -960 420 -950
rect 40 -970 390 -960
rect -60 -1060 -20 -1050
rect -60 -1070 -50 -1060
rect -115 -1080 -50 -1070
rect -30 -1080 -20 -1060
rect -115 -1090 -20 -1080
rect -60 -1125 -20 -1115
rect -60 -1145 -50 -1125
rect -30 -1145 -20 -1125
rect -60 -1170 -20 -1145
rect -110 -1180 -20 -1170
rect -110 -1750 -100 -1180
rect -80 -1750 -50 -1180
rect -30 -1750 -20 -1180
rect -110 -1760 -20 -1750
rect 40 -1180 80 -970
rect 380 -980 390 -970
rect 410 -980 420 -960
rect 380 -990 420 -980
rect 135 -1000 185 -990
rect 135 -1030 145 -1000
rect 175 -1030 185 -1000
rect 135 -1040 185 -1030
rect 40 -1750 50 -1180
rect 70 -1750 80 -1180
rect 40 -1760 80 -1750
rect 140 -1180 180 -1040
rect 140 -1750 150 -1180
rect 170 -1750 180 -1180
rect -115 -1810 -25 -1800
rect -115 -1820 -55 -1810
rect -65 -1830 -55 -1820
rect -35 -1830 -25 -1810
rect -65 -1840 -25 -1830
rect 140 -1820 180 -1750
rect 240 -1180 280 -1170
rect 240 -1750 250 -1180
rect 270 -1750 280 -1180
rect 240 -1760 280 -1750
rect 340 -1180 380 -1170
rect 340 -1750 350 -1180
rect 370 -1750 380 -1180
rect 340 -1780 380 -1750
rect 440 -1180 480 -935
rect 500 -960 880 -950
rect 500 -980 510 -960
rect 530 -970 880 -960
rect 530 -980 540 -970
rect 500 -990 540 -980
rect 440 -1750 450 -1180
rect 470 -1750 480 -1180
rect 440 -1760 480 -1750
rect 540 -1035 590 -1025
rect 540 -1065 550 -1035
rect 580 -1065 590 -1035
rect 540 -1075 590 -1065
rect 540 -1180 580 -1075
rect 540 -1750 550 -1180
rect 570 -1750 580 -1180
rect 540 -1780 580 -1750
rect 640 -1180 680 -1170
rect 640 -1750 650 -1180
rect 670 -1750 680 -1180
rect 640 -1760 680 -1750
rect 740 -1180 780 -1170
rect 740 -1750 750 -1180
rect 770 -1750 780 -1180
rect 340 -1800 580 -1780
rect 740 -1820 780 -1750
rect 840 -1180 880 -970
rect 840 -1750 850 -1180
rect 870 -1750 880 -1180
rect 840 -1760 880 -1750
rect 940 -1125 980 -1115
rect 940 -1145 950 -1125
rect 970 -1145 980 -1125
rect 940 -1170 980 -1145
rect 940 -1180 1030 -1170
rect 940 -1750 950 -1180
rect 970 -1750 1000 -1180
rect 1020 -1750 1030 -1180
rect 940 -1760 1030 -1750
rect 140 -1840 780 -1820
<< viali >>
rect -100 -1750 -80 -1180
rect -50 -1750 -30 -1180
rect 145 -1030 175 -1000
rect 250 -1750 270 -1180
rect 550 -1065 580 -1035
rect 650 -1750 670 -1180
rect 950 -1750 970 -1180
rect 1000 -1750 1020 -1180
<< metal1 >>
rect 135 -1000 185 -990
rect 135 -1030 145 -1000
rect 175 -1030 185 -1000
rect 135 -1040 185 -1030
rect 540 -1035 590 -1030
rect 540 -1065 550 -1035
rect 580 -1065 590 -1035
rect 540 -1075 590 -1065
rect -115 -1180 1035 -1170
rect -115 -1750 -100 -1180
rect -80 -1750 -50 -1180
rect -30 -1750 250 -1180
rect 270 -1750 650 -1180
rect 670 -1750 950 -1180
rect 970 -1750 1000 -1180
rect 1020 -1750 1035 -1180
rect -115 -1760 1035 -1750
<< via1 >>
rect 145 -1030 175 -1000
rect 550 -1065 580 -1035
<< metal2 >>
rect 135 -1000 185 -935
rect 135 -1030 145 -1000
rect 175 -1030 185 -1000
rect 135 -1040 185 -1030
rect 540 -1035 590 -935
rect 540 -1065 550 -1035
rect 580 -1065 590 -1035
rect 540 -1075 590 -1065
<< labels >>
rlabel locali -115 -1080 -115 -1080 7 Vcn
rlabel locali -115 -1810 -115 -1810 7 Vbn
rlabel metal1 -115 -1470 -115 -1470 7 Vn
<< end >>
