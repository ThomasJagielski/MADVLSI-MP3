magic
tech sky130A
timestamp 1615655827
<< nwell >>
rect -120 -910 1230 625
<< nmos >>
rect 0 -1750 50 -1150
rect 100 -1750 150 -1150
rect 200 -1750 250 -1150
rect 300 -1750 350 -1150
rect 480 -1750 530 -1150
rect 580 -1750 630 -1150
rect 760 -1750 810 -1150
rect 860 -1750 910 -1150
rect 960 -1750 1010 -1150
rect 1060 -1750 1110 -1150
rect 0 -2630 50 -2030
rect 100 -2630 150 -2030
rect 200 -2630 250 -2030
rect 300 -2630 350 -2030
rect 480 -2630 530 -2030
rect 580 -2630 630 -2030
rect 760 -2630 810 -2030
rect 860 -2630 910 -2030
rect 960 -2630 1010 -2030
rect 1060 -2630 1110 -2030
<< pmos >>
rect 0 0 50 600
rect 100 0 150 600
rect 200 0 250 600
rect 380 0 430 600
rect 480 0 530 600
rect 580 0 630 600
rect 680 0 730 600
rect 860 0 910 600
rect 960 0 1010 600
rect 1060 0 1110 600
rect 0 -885 50 -285
rect 100 -885 150 -285
rect 200 -885 250 -285
rect 300 -885 350 -285
rect 480 -885 530 -285
rect 580 -885 630 -285
rect 760 -885 810 -285
rect 860 -885 910 -285
rect 960 -885 1010 -285
rect 1060 -885 1110 -285
<< ndiff >>
rect -50 -1165 0 -1150
rect -50 -1735 -35 -1165
rect -15 -1735 0 -1165
rect -50 -1750 0 -1735
rect 50 -1165 100 -1150
rect 50 -1735 65 -1165
rect 85 -1735 100 -1165
rect 50 -1750 100 -1735
rect 150 -1165 200 -1150
rect 150 -1735 165 -1165
rect 185 -1735 200 -1165
rect 150 -1750 200 -1735
rect 250 -1165 300 -1150
rect 250 -1735 265 -1165
rect 285 -1735 300 -1165
rect 250 -1750 300 -1735
rect 350 -1165 400 -1150
rect 350 -1735 365 -1165
rect 385 -1735 400 -1165
rect 350 -1750 400 -1735
rect 430 -1165 480 -1150
rect 430 -1735 445 -1165
rect 465 -1735 480 -1165
rect 430 -1750 480 -1735
rect 530 -1165 580 -1150
rect 530 -1735 545 -1165
rect 565 -1735 580 -1165
rect 530 -1750 580 -1735
rect 630 -1165 680 -1150
rect 630 -1735 645 -1165
rect 665 -1735 680 -1165
rect 630 -1750 680 -1735
rect 710 -1165 760 -1150
rect 710 -1735 725 -1165
rect 745 -1735 760 -1165
rect 710 -1750 760 -1735
rect 810 -1165 860 -1150
rect 810 -1735 825 -1165
rect 845 -1735 860 -1165
rect 810 -1750 860 -1735
rect 910 -1165 960 -1150
rect 910 -1735 925 -1165
rect 945 -1735 960 -1165
rect 910 -1750 960 -1735
rect 1010 -1165 1060 -1150
rect 1010 -1735 1025 -1165
rect 1045 -1735 1060 -1165
rect 1010 -1750 1060 -1735
rect 1110 -1165 1160 -1150
rect 1110 -1735 1125 -1165
rect 1145 -1735 1160 -1165
rect 1110 -1750 1160 -1735
rect -50 -2045 0 -2030
rect -50 -2615 -35 -2045
rect -15 -2615 0 -2045
rect -50 -2630 0 -2615
rect 50 -2045 100 -2030
rect 50 -2615 65 -2045
rect 85 -2615 100 -2045
rect 50 -2630 100 -2615
rect 150 -2045 200 -2030
rect 150 -2615 165 -2045
rect 185 -2615 200 -2045
rect 150 -2630 200 -2615
rect 250 -2045 300 -2030
rect 250 -2615 265 -2045
rect 285 -2615 300 -2045
rect 250 -2630 300 -2615
rect 350 -2045 400 -2030
rect 350 -2615 365 -2045
rect 385 -2615 400 -2045
rect 350 -2630 400 -2615
rect 430 -2045 480 -2030
rect 430 -2615 445 -2045
rect 465 -2615 480 -2045
rect 430 -2630 480 -2615
rect 530 -2045 580 -2030
rect 530 -2615 545 -2045
rect 565 -2615 580 -2045
rect 530 -2630 580 -2615
rect 630 -2045 680 -2030
rect 630 -2615 645 -2045
rect 665 -2615 680 -2045
rect 630 -2630 680 -2615
rect 710 -2045 760 -2030
rect 710 -2615 725 -2045
rect 745 -2615 760 -2045
rect 710 -2630 760 -2615
rect 810 -2045 860 -2030
rect 810 -2615 825 -2045
rect 845 -2615 860 -2045
rect 810 -2630 860 -2615
rect 910 -2045 960 -2030
rect 910 -2615 925 -2045
rect 945 -2615 960 -2045
rect 910 -2630 960 -2615
rect 1010 -2045 1060 -2030
rect 1010 -2615 1025 -2045
rect 1045 -2615 1060 -2045
rect 1010 -2630 1060 -2615
rect 1110 -2045 1160 -2030
rect 1110 -2615 1125 -2045
rect 1145 -2615 1160 -2045
rect 1110 -2630 1160 -2615
<< pdiff >>
rect -50 585 0 600
rect -50 15 -35 585
rect -15 15 0 585
rect -50 0 0 15
rect 50 585 100 600
rect 50 15 65 585
rect 85 15 100 585
rect 50 0 100 15
rect 150 585 200 600
rect 150 15 165 585
rect 185 15 200 585
rect 150 0 200 15
rect 250 585 300 600
rect 250 15 265 585
rect 285 15 300 585
rect 250 0 300 15
rect 330 585 380 600
rect 330 15 345 585
rect 365 15 380 585
rect 330 0 380 15
rect 430 585 480 600
rect 430 15 445 585
rect 465 15 480 585
rect 430 0 480 15
rect 530 585 580 600
rect 530 15 545 585
rect 565 15 580 585
rect 530 0 580 15
rect 630 585 680 600
rect 630 15 645 585
rect 665 15 680 585
rect 630 0 680 15
rect 730 585 780 600
rect 730 15 745 585
rect 765 15 780 585
rect 730 0 780 15
rect 810 585 860 600
rect 810 15 825 585
rect 845 15 860 585
rect 810 0 860 15
rect 910 585 960 600
rect 910 15 925 585
rect 945 15 960 585
rect 910 0 960 15
rect 1010 585 1060 600
rect 1010 15 1025 585
rect 1045 15 1060 585
rect 1010 0 1060 15
rect 1110 585 1160 600
rect 1110 15 1125 585
rect 1145 15 1160 585
rect 1110 0 1160 15
rect -50 -300 0 -285
rect -50 -870 -35 -300
rect -15 -870 0 -300
rect -50 -885 0 -870
rect 50 -300 100 -285
rect 50 -870 65 -300
rect 85 -870 100 -300
rect 50 -885 100 -870
rect 150 -300 200 -285
rect 150 -870 165 -300
rect 185 -870 200 -300
rect 150 -885 200 -870
rect 250 -300 300 -285
rect 250 -870 265 -300
rect 285 -870 300 -300
rect 250 -885 300 -870
rect 350 -300 400 -285
rect 350 -870 365 -300
rect 385 -870 400 -300
rect 350 -885 400 -870
rect 430 -300 480 -285
rect 430 -870 445 -300
rect 465 -870 480 -300
rect 430 -885 480 -870
rect 530 -300 580 -285
rect 530 -870 545 -300
rect 565 -870 580 -300
rect 530 -885 580 -870
rect 630 -300 680 -285
rect 630 -870 645 -300
rect 665 -870 680 -300
rect 630 -885 680 -870
rect 710 -300 760 -285
rect 710 -870 725 -300
rect 745 -870 760 -300
rect 710 -885 760 -870
rect 810 -300 860 -285
rect 810 -870 825 -300
rect 845 -870 860 -300
rect 810 -885 860 -870
rect 910 -300 960 -285
rect 910 -870 925 -300
rect 945 -870 960 -300
rect 910 -885 960 -870
rect 1010 -300 1060 -285
rect 1010 -870 1025 -300
rect 1045 -870 1060 -300
rect 1010 -885 1060 -870
rect 1110 -300 1160 -285
rect 1110 -870 1125 -300
rect 1145 -870 1160 -300
rect 1110 -885 1160 -870
<< ndiffc >>
rect -35 -1735 -15 -1165
rect 65 -1735 85 -1165
rect 165 -1735 185 -1165
rect 265 -1735 285 -1165
rect 365 -1735 385 -1165
rect 445 -1735 465 -1165
rect 545 -1735 565 -1165
rect 645 -1735 665 -1165
rect 725 -1735 745 -1165
rect 825 -1735 845 -1165
rect 925 -1735 945 -1165
rect 1025 -1735 1045 -1165
rect 1125 -1735 1145 -1165
rect -35 -2615 -15 -2045
rect 65 -2615 85 -2045
rect 165 -2615 185 -2045
rect 265 -2615 285 -2045
rect 365 -2615 385 -2045
rect 445 -2615 465 -2045
rect 545 -2615 565 -2045
rect 645 -2615 665 -2045
rect 725 -2615 745 -2045
rect 825 -2615 845 -2045
rect 925 -2615 945 -2045
rect 1025 -2615 1045 -2045
rect 1125 -2615 1145 -2045
<< pdiffc >>
rect -35 15 -15 585
rect 65 15 85 585
rect 165 15 185 585
rect 265 15 285 585
rect 345 15 365 585
rect 445 15 465 585
rect 545 15 565 585
rect 645 15 665 585
rect 745 15 765 585
rect 825 15 845 585
rect 925 15 945 585
rect 1025 15 1045 585
rect 1125 15 1145 585
rect -35 -870 -15 -300
rect 65 -870 85 -300
rect 165 -870 185 -300
rect 265 -870 285 -300
rect 365 -870 385 -300
rect 445 -870 465 -300
rect 545 -870 565 -300
rect 645 -870 665 -300
rect 725 -870 745 -300
rect 825 -870 845 -300
rect 925 -870 945 -300
rect 1025 -870 1045 -300
rect 1125 -870 1145 -300
<< psubdiff >>
rect -100 -1165 -50 -1150
rect -100 -1735 -85 -1165
rect -65 -1735 -50 -1165
rect -100 -1750 -50 -1735
rect 1160 -1165 1210 -1150
rect 1160 -1735 1175 -1165
rect 1195 -1735 1210 -1165
rect 1160 -1750 1210 -1735
rect -100 -2045 -50 -2030
rect -100 -2615 -85 -2045
rect -65 -2615 -50 -2045
rect -100 -2630 -50 -2615
rect 1160 -2045 1210 -2030
rect 1160 -2615 1175 -2045
rect 1195 -2615 1210 -2045
rect 1160 -2630 1210 -2615
<< nsubdiff >>
rect -100 585 -50 600
rect -100 15 -85 585
rect -65 15 -50 585
rect -100 0 -50 15
rect 1160 585 1210 600
rect 1160 15 1175 585
rect 1195 15 1210 585
rect 1160 0 1210 15
rect -100 -300 -50 -285
rect -100 -870 -85 -300
rect -65 -870 -50 -300
rect -100 -885 -50 -870
rect 1160 -300 1210 -285
rect 1160 -870 1175 -300
rect 1195 -870 1210 -300
rect 1160 -885 1210 -870
<< psubdiffcont >>
rect -85 -1735 -65 -1165
rect 1175 -1735 1195 -1165
rect -85 -2615 -65 -2045
rect 1175 -2615 1195 -2045
<< nsubdiffcont >>
rect -85 15 -65 585
rect 1175 15 1195 585
rect -85 -870 -65 -300
rect 1175 -870 1195 -300
<< poly >>
rect 0 600 50 615
rect 100 600 150 615
rect 200 600 250 615
rect 380 600 430 615
rect 480 600 530 615
rect 580 600 630 615
rect 680 600 730 615
rect 860 600 910 615
rect 960 600 1010 615
rect 1060 600 1110 615
rect 0 -15 50 0
rect -50 -25 50 -15
rect -50 -45 -40 -25
rect -20 -45 50 -25
rect -50 -55 50 -45
rect 100 -10 150 0
rect 200 -10 250 0
rect 380 -10 430 0
rect 480 -10 530 0
rect 580 -10 630 0
rect 680 -10 730 0
rect 860 -10 910 0
rect 960 -10 1010 0
rect 100 -25 1010 -10
rect 100 -80 115 -25
rect -50 -90 115 -80
rect -50 -110 -40 -90
rect -20 -95 115 -90
rect 995 -85 1010 -25
rect 1060 -15 1110 0
rect 1060 -30 1160 -15
rect 1060 -50 1130 -30
rect 1150 -50 1160 -30
rect 1060 -60 1160 -50
rect 995 -95 1160 -85
rect -20 -110 -10 -95
rect 995 -100 1130 -95
rect -50 -120 -10 -110
rect 1120 -115 1130 -100
rect 1150 -115 1160 -95
rect 1120 -125 1160 -115
rect 55 -240 95 -230
rect 55 -260 65 -240
rect 85 -260 95 -240
rect 355 -240 395 -230
rect 355 -255 365 -240
rect 200 -260 365 -255
rect 385 -260 395 -240
rect 535 -240 575 -230
rect 535 -260 545 -240
rect 565 -260 575 -240
rect 715 -240 755 -230
rect 715 -260 725 -240
rect 745 -255 755 -240
rect 1015 -240 1055 -230
rect 745 -260 910 -255
rect 1015 -260 1025 -240
rect 1045 -260 1055 -240
rect 0 -275 150 -260
rect 0 -285 50 -275
rect 100 -285 150 -275
rect 200 -270 395 -260
rect 200 -285 250 -270
rect 300 -285 350 -270
rect 480 -275 630 -260
rect 715 -270 910 -260
rect 480 -285 530 -275
rect 580 -285 630 -275
rect 760 -285 810 -270
rect 860 -285 910 -270
rect 960 -275 1110 -260
rect 960 -285 1010 -275
rect 1060 -285 1110 -275
rect 0 -900 50 -885
rect 100 -900 150 -885
rect 200 -1045 250 -885
rect 300 -900 350 -885
rect 480 -900 530 -885
rect 580 -950 630 -885
rect 760 -900 810 -885
rect 860 -900 910 -885
rect 960 -900 1010 -885
rect 1060 -900 1110 -885
rect 580 -970 595 -950
rect 615 -970 630 -950
rect 580 -980 630 -970
rect 860 -1005 950 -995
rect 860 -1025 920 -1005
rect 940 -1025 950 -1005
rect 860 -1035 950 -1025
rect 200 -1065 215 -1045
rect 235 -1065 250 -1045
rect 200 -1075 250 -1065
rect 475 -1045 515 -1035
rect 475 -1065 485 -1045
rect 505 -1060 515 -1045
rect 595 -1045 635 -1035
rect 595 -1060 605 -1045
rect 505 -1065 605 -1060
rect 625 -1065 635 -1045
rect 475 -1075 635 -1065
rect 55 -1105 95 -1095
rect 55 -1120 65 -1105
rect 0 -1125 65 -1120
rect 85 -1120 95 -1105
rect 355 -1105 395 -1095
rect 355 -1120 365 -1105
rect 85 -1125 150 -1120
rect 0 -1135 150 -1125
rect 0 -1150 50 -1135
rect 100 -1150 150 -1135
rect 200 -1125 365 -1120
rect 385 -1120 395 -1105
rect 715 -1105 755 -1095
rect 715 -1120 725 -1105
rect 385 -1125 725 -1120
rect 745 -1120 755 -1105
rect 860 -1120 910 -1035
rect 1015 -1105 1055 -1095
rect 1015 -1120 1025 -1105
rect 745 -1125 910 -1120
rect 200 -1135 910 -1125
rect 200 -1150 250 -1135
rect 300 -1150 350 -1135
rect 480 -1150 530 -1135
rect 580 -1150 630 -1135
rect 760 -1150 810 -1135
rect 860 -1150 910 -1135
rect 960 -1125 1025 -1120
rect 1045 -1120 1055 -1105
rect 1045 -1125 1110 -1120
rect 960 -1135 1110 -1125
rect 960 -1150 1010 -1135
rect 1060 -1150 1110 -1135
rect 0 -1765 50 -1750
rect 100 -1765 150 -1750
rect 200 -1765 250 -1750
rect 300 -1765 350 -1750
rect 480 -1765 530 -1750
rect 580 -1765 630 -1750
rect 760 -1765 810 -1750
rect 860 -1765 910 -1750
rect 960 -1765 1010 -1750
rect 1060 -1765 1110 -1750
rect 335 -1975 395 -1965
rect 55 -1985 95 -1975
rect 55 -2000 65 -1985
rect 0 -2005 65 -2000
rect 85 -2000 95 -1985
rect 335 -1995 365 -1975
rect 385 -1985 755 -1975
rect 385 -1990 725 -1985
rect 385 -1995 395 -1990
rect 335 -2000 395 -1995
rect 85 -2005 150 -2000
rect 0 -2015 150 -2005
rect 0 -2030 50 -2015
rect 100 -2030 150 -2015
rect 200 -2005 395 -2000
rect 715 -2005 725 -1990
rect 745 -2000 755 -1985
rect 1015 -1985 1055 -1975
rect 1015 -2000 1025 -1985
rect 745 -2005 910 -2000
rect 200 -2015 350 -2005
rect 715 -2015 910 -2005
rect 200 -2030 250 -2015
rect 300 -2030 350 -2015
rect 480 -2030 530 -2015
rect 580 -2030 630 -2015
rect 760 -2030 810 -2015
rect 860 -2030 910 -2015
rect 960 -2005 1025 -2000
rect 1045 -2000 1055 -1985
rect 1045 -2005 1110 -2000
rect 960 -2015 1110 -2005
rect 960 -2030 1010 -2015
rect 1060 -2030 1110 -2015
rect 0 -2645 50 -2630
rect 100 -2645 150 -2630
rect 200 -2645 250 -2630
rect 300 -2645 350 -2630
rect 480 -2645 530 -2630
rect 580 -2645 630 -2630
rect 760 -2645 810 -2630
rect 860 -2645 910 -2630
rect 960 -2645 1010 -2630
rect 1060 -2645 1110 -2630
rect 480 -2655 630 -2645
rect 480 -2665 545 -2655
rect 535 -2675 545 -2665
rect 565 -2665 630 -2655
rect 565 -2675 575 -2665
rect 535 -2685 575 -2675
<< polycont >>
rect -40 -45 -20 -25
rect -40 -110 -20 -90
rect 1130 -50 1150 -30
rect 1130 -115 1150 -95
rect 65 -260 85 -240
rect 365 -260 385 -240
rect 545 -260 565 -240
rect 725 -260 745 -240
rect 1025 -260 1045 -240
rect 595 -970 615 -950
rect 920 -1025 940 -1005
rect 215 -1065 235 -1045
rect 485 -1065 505 -1045
rect 605 -1065 625 -1045
rect 65 -1125 85 -1105
rect 365 -1125 385 -1105
rect 725 -1125 745 -1105
rect 1025 -1125 1045 -1105
rect 65 -2005 85 -1985
rect 365 -1995 385 -1975
rect 725 -2005 745 -1985
rect 1025 -2005 1045 -1985
rect 545 -2675 565 -2655
<< locali >>
rect -95 585 -5 595
rect -95 15 -85 585
rect -65 15 -35 585
rect -15 15 -5 585
rect -95 5 -5 15
rect -50 -25 -5 5
rect -50 -45 -40 -25
rect -20 -45 -5 -25
rect -50 -55 -5 -45
rect 55 585 95 595
rect 55 15 65 585
rect 85 15 95 585
rect 55 -80 95 15
rect 155 585 195 595
rect 155 15 165 585
rect 185 15 195 585
rect 155 5 195 15
rect 255 585 295 595
rect 255 15 265 585
rect 285 15 295 585
rect -100 -90 95 -80
rect -100 -110 -40 -90
rect -20 -100 95 -90
rect -20 -110 -10 -100
rect -100 -120 -10 -110
rect 255 -140 295 15
rect 335 585 375 595
rect 335 15 345 585
rect 365 15 375 585
rect 335 -110 375 15
rect 435 585 475 595
rect 435 15 445 585
rect 465 15 475 585
rect 435 10 475 15
rect 535 585 575 595
rect 535 15 545 585
rect 565 15 575 585
rect 535 -60 575 15
rect 635 585 675 595
rect 635 15 645 585
rect 665 15 675 585
rect 635 10 675 15
rect 735 585 775 595
rect 735 15 745 585
rect 765 15 775 585
rect 535 -80 545 -60
rect 565 -80 575 -60
rect 535 -90 575 -80
rect 735 -100 775 15
rect 735 -110 745 -100
rect 335 -120 745 -110
rect 765 -120 775 -100
rect 335 -130 775 -120
rect 815 585 855 595
rect 815 15 825 585
rect 845 15 855 585
rect 255 -160 265 -140
rect 285 -150 295 -140
rect 815 -150 855 15
rect 915 585 955 595
rect 915 15 925 585
rect 945 15 955 585
rect 915 5 955 15
rect 1015 585 1055 595
rect 1015 15 1025 585
rect 1045 15 1055 585
rect 1015 -85 1055 15
rect 1115 585 1205 595
rect 1115 15 1125 585
rect 1145 15 1175 585
rect 1195 15 1205 585
rect 1115 5 1205 15
rect 1115 -30 1160 5
rect 1115 -50 1130 -30
rect 1150 -50 1160 -30
rect 1115 -60 1160 -50
rect 1015 -95 1210 -85
rect 1015 -105 1130 -95
rect 1120 -115 1130 -105
rect 1150 -115 1210 -95
rect 1120 -125 1210 -115
rect 285 -160 855 -150
rect 255 -170 855 -160
rect 355 -210 755 -190
rect -50 -240 95 -230
rect -50 -250 65 -240
rect -50 -290 -5 -250
rect -95 -300 -5 -290
rect -95 -870 -85 -300
rect -65 -870 -35 -300
rect -15 -870 -5 -300
rect -95 -880 -5 -870
rect 55 -260 65 -250
rect 85 -260 95 -240
rect 55 -300 95 -260
rect 355 -240 395 -210
rect 355 -260 365 -240
rect 385 -260 395 -240
rect 55 -870 65 -300
rect 85 -870 95 -300
rect 55 -880 95 -870
rect 155 -300 195 -290
rect 155 -870 165 -300
rect 185 -870 195 -300
rect 155 -880 195 -870
rect 255 -300 295 -290
rect 255 -870 265 -300
rect 285 -870 295 -300
rect 255 -900 295 -870
rect 355 -300 395 -260
rect 535 -240 575 -230
rect 535 -260 545 -240
rect 565 -260 575 -240
rect 355 -870 365 -300
rect 385 -870 395 -300
rect 355 -880 395 -870
rect 435 -300 475 -290
rect 435 -870 445 -300
rect 465 -870 475 -300
rect 435 -900 475 -870
rect 535 -300 575 -260
rect 715 -240 755 -210
rect 715 -260 725 -240
rect 745 -260 755 -240
rect 535 -870 545 -300
rect 565 -870 575 -300
rect 535 -880 575 -870
rect 635 -300 675 -290
rect 635 -870 645 -300
rect 665 -870 675 -300
rect 635 -900 675 -870
rect 715 -300 755 -260
rect 1015 -240 1160 -230
rect 1015 -260 1025 -240
rect 1045 -250 1160 -240
rect 1045 -260 1055 -250
rect 715 -870 725 -300
rect 745 -870 755 -300
rect 715 -880 755 -870
rect 815 -300 855 -290
rect 815 -870 825 -300
rect 845 -870 855 -300
rect 815 -900 855 -870
rect 915 -300 955 -290
rect 915 -870 925 -300
rect 945 -870 955 -300
rect 915 -880 955 -870
rect 1015 -300 1055 -260
rect 1015 -870 1025 -300
rect 1045 -870 1055 -300
rect 1015 -880 1055 -870
rect 1115 -290 1160 -250
rect 1115 -300 1205 -290
rect 1115 -870 1125 -300
rect 1145 -870 1175 -300
rect 1195 -870 1205 -300
rect 1115 -880 1205 -870
rect 255 -920 855 -900
rect 535 -950 1210 -940
rect 535 -970 595 -950
rect 615 -960 1210 -950
rect 615 -970 630 -960
rect 535 -980 630 -970
rect 200 -1045 250 -1035
rect 200 -1055 215 -1045
rect 155 -1065 215 -1055
rect 235 -1055 250 -1045
rect 475 -1045 515 -1035
rect 475 -1055 485 -1045
rect 235 -1065 485 -1055
rect 505 -1065 515 -1045
rect 155 -1075 515 -1065
rect -50 -1105 95 -1095
rect -50 -1115 65 -1105
rect -50 -1155 -5 -1115
rect -95 -1165 -5 -1155
rect -95 -1735 -85 -1165
rect -65 -1735 -35 -1165
rect -15 -1735 -5 -1165
rect -95 -1745 -5 -1735
rect 55 -1125 65 -1115
rect 85 -1125 95 -1105
rect 55 -1165 95 -1125
rect 55 -1735 65 -1165
rect 85 -1735 95 -1165
rect 55 -1745 95 -1735
rect 155 -1165 195 -1075
rect 355 -1105 395 -1095
rect 355 -1125 365 -1105
rect 385 -1125 395 -1105
rect 155 -1735 165 -1165
rect 185 -1735 195 -1165
rect 155 -1745 195 -1735
rect 255 -1165 295 -1155
rect 255 -1735 265 -1165
rect 285 -1735 295 -1165
rect 255 -1765 295 -1735
rect 355 -1165 395 -1125
rect 355 -1735 365 -1165
rect 385 -1735 395 -1165
rect 355 -1745 395 -1735
rect 435 -1165 475 -1155
rect 435 -1735 445 -1165
rect 465 -1735 475 -1165
rect 435 -1765 475 -1735
rect 535 -1165 575 -980
rect 910 -1005 950 -995
rect 910 -1025 920 -1005
rect 940 -1015 950 -1005
rect 940 -1025 1210 -1015
rect 910 -1035 1210 -1025
rect 595 -1045 635 -1035
rect 595 -1065 605 -1045
rect 625 -1055 635 -1045
rect 625 -1065 955 -1055
rect 595 -1075 955 -1065
rect 715 -1105 755 -1095
rect 715 -1125 725 -1105
rect 745 -1125 755 -1105
rect 535 -1735 545 -1165
rect 565 -1735 575 -1165
rect 535 -1745 575 -1735
rect 635 -1165 675 -1155
rect 635 -1735 645 -1165
rect 665 -1735 675 -1165
rect 635 -1765 675 -1735
rect 715 -1165 755 -1125
rect 715 -1735 725 -1165
rect 745 -1735 755 -1165
rect 715 -1745 755 -1735
rect 815 -1165 855 -1155
rect 815 -1735 825 -1165
rect 845 -1735 855 -1165
rect 815 -1765 855 -1735
rect 915 -1165 955 -1075
rect 915 -1735 925 -1165
rect 945 -1735 955 -1165
rect 915 -1745 955 -1735
rect 1015 -1105 1160 -1095
rect 1015 -1125 1025 -1105
rect 1045 -1115 1160 -1105
rect 1045 -1125 1055 -1115
rect 1015 -1165 1055 -1125
rect 1015 -1735 1025 -1165
rect 1045 -1735 1055 -1165
rect 1015 -1745 1055 -1735
rect 1115 -1155 1160 -1115
rect 1115 -1165 1205 -1155
rect 1115 -1735 1125 -1165
rect 1145 -1735 1175 -1165
rect 1195 -1735 1205 -1165
rect 1115 -1745 1205 -1735
rect 255 -1805 855 -1765
rect 255 -1900 855 -1880
rect -50 -1985 95 -1975
rect -50 -1995 65 -1985
rect -50 -2035 -5 -1995
rect 55 -2005 65 -1995
rect 85 -2005 95 -1985
rect 55 -2015 95 -2005
rect -95 -2045 -5 -2035
rect -95 -2615 -85 -2045
rect -65 -2615 -35 -2045
rect -15 -2615 -5 -2045
rect -95 -2625 -5 -2615
rect 55 -2045 95 -2035
rect 55 -2615 65 -2045
rect 85 -2615 95 -2045
rect 55 -2625 95 -2615
rect 155 -2045 195 -2035
rect 155 -2615 165 -2045
rect 185 -2615 195 -2045
rect 155 -2625 195 -2615
rect 255 -2045 295 -1900
rect 255 -2615 265 -2045
rect 285 -2615 295 -2045
rect 255 -2625 295 -2615
rect 355 -1975 395 -1965
rect 355 -1995 365 -1975
rect 385 -1995 395 -1975
rect 355 -2045 395 -1995
rect 355 -2615 365 -2045
rect 385 -2615 395 -2045
rect 355 -2625 395 -2615
rect 435 -2045 475 -1900
rect 435 -2615 445 -2045
rect 465 -2615 475 -2045
rect 435 -2625 475 -2615
rect 535 -1930 575 -1920
rect 535 -1950 545 -1930
rect 565 -1950 575 -1930
rect 535 -2045 575 -1950
rect 535 -2615 545 -2045
rect 565 -2615 575 -2045
rect 535 -2655 575 -2615
rect 635 -2045 675 -1900
rect 635 -2615 645 -2045
rect 665 -2615 675 -2045
rect 635 -2625 675 -2615
rect 715 -1985 755 -1975
rect 715 -2005 725 -1985
rect 745 -2005 755 -1985
rect 715 -2045 755 -2005
rect 715 -2615 725 -2045
rect 745 -2615 755 -2045
rect 715 -2625 755 -2615
rect 815 -2045 855 -1900
rect 1015 -1985 1160 -1975
rect 1015 -2005 1025 -1985
rect 1045 -2000 1160 -1985
rect 1045 -2005 1055 -2000
rect 815 -2615 825 -2045
rect 845 -2615 855 -2045
rect 815 -2625 855 -2615
rect 915 -2045 955 -2035
rect 915 -2615 925 -2045
rect 945 -2615 955 -2045
rect 915 -2625 955 -2615
rect 1015 -2045 1055 -2005
rect 1015 -2615 1025 -2045
rect 1045 -2615 1055 -2045
rect 1015 -2625 1055 -2615
rect 1115 -2035 1160 -2000
rect 1115 -2045 1205 -2035
rect 1115 -2615 1125 -2045
rect 1145 -2615 1175 -2045
rect 1195 -2615 1205 -2045
rect 1115 -2625 1205 -2615
rect 535 -2675 545 -2655
rect 565 -2665 575 -2655
rect 565 -2675 1210 -2665
rect 535 -2685 1210 -2675
<< viali >>
rect -85 15 -65 585
rect -35 15 -15 585
rect 165 15 185 585
rect 445 15 465 585
rect 645 15 665 585
rect 545 -80 565 -60
rect 745 -120 765 -100
rect 265 -160 285 -140
rect 925 15 945 585
rect 1125 15 1145 585
rect 1175 15 1195 585
rect -85 -870 -65 -300
rect -35 -870 -15 -300
rect 65 -870 85 -300
rect 165 -870 185 -300
rect 925 -870 945 -300
rect 1025 -870 1045 -300
rect 1125 -870 1145 -300
rect 1175 -870 1195 -300
rect -85 -1735 -65 -1165
rect -35 -1735 -15 -1165
rect 65 -1735 85 -1165
rect 365 -1125 385 -1105
rect 265 -1735 285 -1165
rect 825 -1735 845 -1165
rect 1025 -1735 1045 -1165
rect 1125 -1735 1145 -1165
rect 1175 -1735 1195 -1165
rect -85 -2615 -65 -2045
rect -35 -2615 -15 -2045
rect 65 -2615 85 -2045
rect 165 -2615 185 -2045
rect 365 -1995 385 -1975
rect 545 -1950 565 -1930
rect 925 -2615 945 -2045
rect 1025 -2615 1045 -2045
rect 1125 -2615 1145 -2045
rect 1175 -2615 1195 -2045
<< metal1 >>
rect -100 585 1210 595
rect -100 15 -85 585
rect -65 15 -35 585
rect -15 15 165 585
rect 185 15 445 585
rect 465 15 645 585
rect 665 15 925 585
rect 945 15 1125 585
rect 1145 15 1175 585
rect 1195 15 1210 585
rect -100 5 1210 15
rect -100 -300 195 5
rect 535 -60 575 -50
rect 535 -80 545 -60
rect 565 -80 575 -60
rect -100 -870 -85 -300
rect -65 -870 -35 -300
rect -15 -870 65 -300
rect 85 -870 165 -300
rect 185 -870 195 -300
rect -100 -880 195 -870
rect 255 -140 295 -130
rect 255 -160 265 -140
rect 285 -160 295 -140
rect 255 -1095 295 -160
rect 255 -1105 395 -1095
rect 255 -1125 365 -1105
rect 385 -1125 395 -1105
rect 355 -1135 395 -1125
rect -100 -1165 300 -1155
rect -100 -1735 -85 -1165
rect -65 -1735 -35 -1165
rect -15 -1735 65 -1165
rect 85 -1735 265 -1165
rect 285 -1735 300 -1165
rect -100 -2035 300 -1735
rect 535 -1765 575 -80
rect 355 -1805 575 -1765
rect 735 -100 775 -90
rect 735 -120 745 -100
rect 765 -120 775 -100
rect 355 -1975 395 -1805
rect 735 -1920 775 -120
rect 915 -300 1210 5
rect 915 -870 925 -300
rect 945 -870 1025 -300
rect 1045 -870 1125 -300
rect 1145 -870 1175 -300
rect 1195 -870 1210 -300
rect 915 -880 1210 -870
rect 535 -1930 775 -1920
rect 535 -1950 545 -1930
rect 565 -1950 775 -1930
rect 535 -1960 775 -1950
rect 810 -1165 1210 -1155
rect 810 -1735 825 -1165
rect 845 -1735 1025 -1165
rect 1045 -1735 1125 -1165
rect 1145 -1735 1175 -1165
rect 1195 -1735 1210 -1165
rect 355 -1995 365 -1975
rect 385 -1995 395 -1975
rect 355 -2005 395 -1995
rect 810 -2035 1210 -1735
rect -100 -2045 1210 -2035
rect -100 -2615 -85 -2045
rect -65 -2615 -35 -2045
rect -15 -2615 65 -2045
rect 85 -2615 165 -2045
rect 185 -2615 925 -2045
rect 945 -2615 1025 -2045
rect 1045 -2615 1125 -2045
rect 1145 -2615 1175 -2045
rect 1195 -2615 1210 -2045
rect -100 -2625 1210 -2615
<< labels >>
rlabel locali -100 -100 -100 -100 7 Vbp
rlabel metal1 -100 300 -100 300 7 VP
rlabel metal1 -100 -2330 -100 -2330 7 VN
rlabel locali 1210 -2675 1210 -2675 3 Vcn
rlabel locali 1210 -950 1210 -950 3 Vcp
rlabel locali 1210 -1025 1210 -1025 3 Vbn
<< end >>
