magic
tech sky130A
timestamp 1615694345
<< nwell >>
rect -120 -935 1230 635
<< nmos >>
rect 0 -1750 50 -1150
rect 100 -1750 150 -1150
rect 200 -1750 250 -1150
rect 300 -1750 350 -1150
rect 480 -1750 530 -1150
rect 580 -1750 630 -1150
rect 760 -1750 810 -1150
rect 860 -1750 910 -1150
rect 960 -1750 1010 -1150
rect 1060 -1750 1110 -1150
rect 0 -2575 50 -1975
rect 100 -2575 150 -1975
rect 200 -2575 250 -1975
rect 300 -2575 350 -1975
rect 480 -2575 530 -1975
rect 580 -2575 630 -1975
rect 760 -2575 810 -1975
rect 860 -2575 910 -1975
rect 960 -2575 1010 -1975
rect 1060 -2575 1110 -1975
<< pmos >>
rect 0 15 50 615
rect 100 15 150 615
rect 200 15 250 615
rect 380 15 430 615
rect 480 15 530 615
rect 580 15 630 615
rect 680 15 730 615
rect 860 15 910 615
rect 960 15 1010 615
rect 1060 15 1110 615
rect 0 -915 50 -315
rect 100 -915 150 -315
rect 200 -915 250 -315
rect 300 -915 350 -315
rect 480 -915 530 -315
rect 580 -915 630 -315
rect 760 -915 810 -315
rect 860 -915 910 -315
rect 960 -915 1010 -315
rect 1060 -915 1110 -315
<< ndiff >>
rect -50 -1165 0 -1150
rect -50 -1735 -35 -1165
rect -15 -1735 0 -1165
rect -50 -1750 0 -1735
rect 50 -1165 100 -1150
rect 50 -1735 65 -1165
rect 85 -1735 100 -1165
rect 50 -1750 100 -1735
rect 150 -1165 200 -1150
rect 150 -1735 165 -1165
rect 185 -1735 200 -1165
rect 150 -1750 200 -1735
rect 250 -1165 300 -1150
rect 250 -1735 265 -1165
rect 285 -1735 300 -1165
rect 250 -1750 300 -1735
rect 350 -1165 400 -1150
rect 350 -1735 365 -1165
rect 385 -1735 400 -1165
rect 350 -1750 400 -1735
rect 430 -1165 480 -1150
rect 430 -1735 445 -1165
rect 465 -1735 480 -1165
rect 430 -1750 480 -1735
rect 530 -1165 580 -1150
rect 530 -1735 545 -1165
rect 565 -1735 580 -1165
rect 530 -1750 580 -1735
rect 630 -1165 680 -1150
rect 630 -1735 645 -1165
rect 665 -1735 680 -1165
rect 630 -1750 680 -1735
rect 710 -1165 760 -1150
rect 710 -1735 725 -1165
rect 745 -1735 760 -1165
rect 710 -1750 760 -1735
rect 810 -1165 860 -1150
rect 810 -1735 825 -1165
rect 845 -1735 860 -1165
rect 810 -1750 860 -1735
rect 910 -1165 960 -1150
rect 910 -1735 925 -1165
rect 945 -1735 960 -1165
rect 910 -1750 960 -1735
rect 1010 -1165 1060 -1150
rect 1010 -1735 1025 -1165
rect 1045 -1735 1060 -1165
rect 1010 -1750 1060 -1735
rect 1110 -1165 1160 -1150
rect 1110 -1735 1125 -1165
rect 1145 -1735 1160 -1165
rect 1110 -1750 1160 -1735
rect -50 -1990 0 -1975
rect -50 -2560 -35 -1990
rect -15 -2560 0 -1990
rect -50 -2575 0 -2560
rect 50 -1990 100 -1975
rect 50 -2560 65 -1990
rect 85 -2560 100 -1990
rect 50 -2575 100 -2560
rect 150 -1990 200 -1975
rect 150 -2560 165 -1990
rect 185 -2560 200 -1990
rect 150 -2575 200 -2560
rect 250 -1990 300 -1975
rect 250 -2560 265 -1990
rect 285 -2560 300 -1990
rect 250 -2575 300 -2560
rect 350 -1990 400 -1975
rect 350 -2560 365 -1990
rect 385 -2560 400 -1990
rect 350 -2575 400 -2560
rect 430 -1990 480 -1975
rect 430 -2560 445 -1990
rect 465 -2560 480 -1990
rect 430 -2575 480 -2560
rect 530 -1990 580 -1975
rect 530 -2560 545 -1990
rect 565 -2560 580 -1990
rect 530 -2575 580 -2560
rect 630 -1990 680 -1975
rect 630 -2560 645 -1990
rect 665 -2560 680 -1990
rect 630 -2575 680 -2560
rect 710 -1990 760 -1975
rect 710 -2560 725 -1990
rect 745 -2560 760 -1990
rect 710 -2575 760 -2560
rect 810 -1990 860 -1975
rect 810 -2560 825 -1990
rect 845 -2560 860 -1990
rect 810 -2575 860 -2560
rect 910 -1990 960 -1975
rect 910 -2560 925 -1990
rect 945 -2560 960 -1990
rect 910 -2575 960 -2560
rect 1010 -1990 1060 -1975
rect 1010 -2560 1025 -1990
rect 1045 -2560 1060 -1990
rect 1010 -2575 1060 -2560
rect 1110 -1990 1160 -1975
rect 1110 -2560 1125 -1990
rect 1145 -2560 1160 -1990
rect 1110 -2575 1160 -2560
<< pdiff >>
rect -50 600 0 615
rect -50 30 -35 600
rect -15 30 0 600
rect -50 15 0 30
rect 50 600 100 615
rect 50 30 65 600
rect 85 30 100 600
rect 50 15 100 30
rect 150 600 200 615
rect 150 30 165 600
rect 185 30 200 600
rect 150 15 200 30
rect 250 600 300 615
rect 250 30 265 600
rect 285 30 300 600
rect 250 15 300 30
rect 330 600 380 615
rect 330 30 345 600
rect 365 30 380 600
rect 330 15 380 30
rect 430 600 480 615
rect 430 30 445 600
rect 465 30 480 600
rect 430 15 480 30
rect 530 600 580 615
rect 530 30 545 600
rect 565 30 580 600
rect 530 15 580 30
rect 630 600 680 615
rect 630 30 645 600
rect 665 30 680 600
rect 630 15 680 30
rect 730 600 780 615
rect 730 30 745 600
rect 765 30 780 600
rect 730 15 780 30
rect 810 600 860 615
rect 810 30 825 600
rect 845 30 860 600
rect 810 15 860 30
rect 910 600 960 615
rect 910 30 925 600
rect 945 30 960 600
rect 910 15 960 30
rect 1010 600 1060 615
rect 1010 30 1025 600
rect 1045 30 1060 600
rect 1010 15 1060 30
rect 1110 600 1160 615
rect 1110 30 1125 600
rect 1145 30 1160 600
rect 1110 15 1160 30
rect -50 -330 0 -315
rect -50 -900 -35 -330
rect -15 -900 0 -330
rect -50 -915 0 -900
rect 50 -330 100 -315
rect 50 -900 65 -330
rect 85 -900 100 -330
rect 50 -915 100 -900
rect 150 -330 200 -315
rect 150 -900 165 -330
rect 185 -900 200 -330
rect 150 -915 200 -900
rect 250 -330 300 -315
rect 250 -900 265 -330
rect 285 -900 300 -330
rect 250 -915 300 -900
rect 350 -330 400 -315
rect 350 -900 365 -330
rect 385 -900 400 -330
rect 350 -915 400 -900
rect 430 -330 480 -315
rect 430 -900 445 -330
rect 465 -900 480 -330
rect 430 -915 480 -900
rect 530 -330 580 -315
rect 530 -900 545 -330
rect 565 -900 580 -330
rect 530 -915 580 -900
rect 630 -330 680 -315
rect 630 -900 645 -330
rect 665 -900 680 -330
rect 630 -915 680 -900
rect 710 -330 760 -315
rect 710 -900 725 -330
rect 745 -900 760 -330
rect 710 -915 760 -900
rect 810 -330 860 -315
rect 810 -900 825 -330
rect 845 -900 860 -330
rect 810 -915 860 -900
rect 910 -330 960 -315
rect 910 -900 925 -330
rect 945 -900 960 -330
rect 910 -915 960 -900
rect 1010 -330 1060 -315
rect 1010 -900 1025 -330
rect 1045 -900 1060 -330
rect 1010 -915 1060 -900
rect 1110 -330 1160 -315
rect 1110 -900 1125 -330
rect 1145 -900 1160 -330
rect 1110 -915 1160 -900
<< ndiffc >>
rect -35 -1735 -15 -1165
rect 65 -1735 85 -1165
rect 165 -1735 185 -1165
rect 265 -1735 285 -1165
rect 365 -1735 385 -1165
rect 445 -1735 465 -1165
rect 545 -1735 565 -1165
rect 645 -1735 665 -1165
rect 725 -1735 745 -1165
rect 825 -1735 845 -1165
rect 925 -1735 945 -1165
rect 1025 -1735 1045 -1165
rect 1125 -1735 1145 -1165
rect -35 -2560 -15 -1990
rect 65 -2560 85 -1990
rect 165 -2560 185 -1990
rect 265 -2560 285 -1990
rect 365 -2560 385 -1990
rect 445 -2560 465 -1990
rect 545 -2560 565 -1990
rect 645 -2560 665 -1990
rect 725 -2560 745 -1990
rect 825 -2560 845 -1990
rect 925 -2560 945 -1990
rect 1025 -2560 1045 -1990
rect 1125 -2560 1145 -1990
<< pdiffc >>
rect -35 30 -15 600
rect 65 30 85 600
rect 165 30 185 600
rect 265 30 285 600
rect 345 30 365 600
rect 445 30 465 600
rect 545 30 565 600
rect 645 30 665 600
rect 745 30 765 600
rect 825 30 845 600
rect 925 30 945 600
rect 1025 30 1045 600
rect 1125 30 1145 600
rect -35 -900 -15 -330
rect 65 -900 85 -330
rect 165 -900 185 -330
rect 265 -900 285 -330
rect 365 -900 385 -330
rect 445 -900 465 -330
rect 545 -900 565 -330
rect 645 -900 665 -330
rect 725 -900 745 -330
rect 825 -900 845 -330
rect 925 -900 945 -330
rect 1025 -900 1045 -330
rect 1125 -900 1145 -330
<< psubdiff >>
rect -100 -1165 -50 -1150
rect -100 -1735 -85 -1165
rect -65 -1735 -50 -1165
rect -100 -1750 -50 -1735
rect 1160 -1165 1210 -1150
rect 1160 -1735 1175 -1165
rect 1195 -1735 1210 -1165
rect 1160 -1750 1210 -1735
rect -100 -1990 -50 -1975
rect -100 -2560 -85 -1990
rect -65 -2560 -50 -1990
rect -100 -2575 -50 -2560
rect 1160 -1990 1210 -1975
rect 1160 -2560 1175 -1990
rect 1195 -2560 1210 -1990
rect 1160 -2575 1210 -2560
<< nsubdiff >>
rect -100 600 -50 615
rect -100 30 -85 600
rect -65 30 -50 600
rect -100 15 -50 30
rect 1160 600 1210 615
rect 1160 30 1175 600
rect 1195 30 1210 600
rect 1160 15 1210 30
rect -100 -330 -50 -315
rect -100 -900 -85 -330
rect -65 -900 -50 -330
rect -100 -915 -50 -900
rect 1160 -330 1210 -315
rect 1160 -900 1175 -330
rect 1195 -900 1210 -330
rect 1160 -915 1210 -900
<< psubdiffcont >>
rect -85 -1735 -65 -1165
rect 1175 -1735 1195 -1165
rect -85 -2560 -65 -1990
rect 1175 -2560 1195 -1990
<< nsubdiffcont >>
rect -85 30 -65 600
rect 1175 30 1195 600
rect -85 -900 -65 -330
rect 1175 -900 1195 -330
<< poly >>
rect 860 660 910 670
rect 860 640 880 660
rect 900 640 910 660
rect 0 615 50 630
rect 100 615 150 630
rect 200 615 250 630
rect 380 615 430 630
rect 480 615 530 630
rect 580 615 630 630
rect 680 615 730 630
rect 860 615 910 640
rect 960 615 1010 630
rect 1060 615 1110 630
rect 0 0 50 15
rect -50 -10 50 0
rect -50 -30 -40 -10
rect -20 -30 50 -10
rect -50 -40 50 -30
rect 100 5 150 15
rect 200 5 250 15
rect 380 5 430 15
rect 480 5 530 15
rect 580 5 630 15
rect 680 5 730 15
rect 860 5 910 15
rect 960 5 1010 15
rect 100 -10 1010 5
rect 1060 0 1110 15
rect 100 -65 115 -10
rect 1060 -15 1160 0
rect 1060 -35 1130 -15
rect 1150 -35 1160 -15
rect 1060 -45 1160 -35
rect -50 -75 115 -65
rect -50 -95 -40 -75
rect -20 -80 115 -75
rect -20 -95 -10 -80
rect -50 -105 -10 -95
rect 55 -270 95 -260
rect 55 -290 65 -270
rect 85 -290 95 -270
rect 355 -270 395 -260
rect 355 -285 365 -270
rect 200 -290 365 -285
rect 385 -290 395 -270
rect 535 -270 575 -260
rect 535 -290 545 -270
rect 565 -290 575 -270
rect 715 -270 755 -260
rect 715 -290 725 -270
rect 745 -285 755 -270
rect 1015 -270 1055 -260
rect 745 -290 910 -285
rect 1015 -290 1025 -270
rect 1045 -290 1055 -270
rect 0 -305 150 -290
rect 0 -315 50 -305
rect 100 -315 150 -305
rect 200 -300 395 -290
rect 200 -315 250 -300
rect 300 -315 350 -300
rect 480 -305 630 -290
rect 715 -300 910 -290
rect 480 -315 530 -305
rect 580 -315 630 -305
rect 760 -315 810 -300
rect 860 -315 910 -300
rect 960 -305 1110 -290
rect 960 -315 1010 -305
rect 1060 -315 1110 -305
rect 0 -930 50 -915
rect 100 -930 150 -915
rect 200 -1045 250 -915
rect 300 -930 350 -915
rect 480 -930 530 -915
rect 580 -980 630 -915
rect 760 -930 810 -915
rect 860 -930 910 -915
rect 960 -930 1010 -915
rect 1060 -930 1110 -915
rect 580 -1000 595 -980
rect 615 -1000 630 -980
rect 580 -1010 630 -1000
rect 200 -1065 215 -1045
rect 235 -1065 250 -1045
rect 200 -1075 250 -1065
rect 475 -1045 515 -1035
rect 475 -1065 485 -1045
rect 505 -1060 515 -1045
rect 595 -1045 635 -1035
rect 595 -1060 605 -1045
rect 505 -1065 605 -1060
rect 625 -1065 635 -1045
rect 1015 -1040 1055 -1030
rect 1015 -1055 1025 -1040
rect 475 -1075 635 -1065
rect 895 -1060 1025 -1055
rect 1045 -1060 1055 -1040
rect 895 -1070 1055 -1060
rect 55 -1105 95 -1095
rect 55 -1120 65 -1105
rect 0 -1125 65 -1120
rect 85 -1120 95 -1105
rect 355 -1105 395 -1095
rect 355 -1120 365 -1105
rect 85 -1125 150 -1120
rect 0 -1135 150 -1125
rect 0 -1150 50 -1135
rect 100 -1150 150 -1135
rect 200 -1125 365 -1120
rect 385 -1120 395 -1105
rect 715 -1105 755 -1095
rect 715 -1120 725 -1105
rect 385 -1125 725 -1120
rect 745 -1120 755 -1105
rect 895 -1120 910 -1070
rect 1015 -1105 1055 -1095
rect 1015 -1120 1025 -1105
rect 745 -1125 910 -1120
rect 200 -1135 910 -1125
rect 200 -1150 250 -1135
rect 300 -1150 350 -1135
rect 480 -1150 530 -1135
rect 580 -1150 630 -1135
rect 760 -1150 810 -1135
rect 860 -1150 910 -1135
rect 960 -1125 1025 -1120
rect 1045 -1120 1055 -1105
rect 1045 -1125 1110 -1120
rect 960 -1135 1110 -1125
rect 960 -1150 1010 -1135
rect 1060 -1150 1110 -1135
rect 0 -1765 50 -1750
rect 100 -1765 150 -1750
rect 200 -1765 250 -1750
rect 300 -1765 350 -1750
rect 480 -1765 530 -1750
rect 580 -1765 630 -1750
rect 760 -1765 810 -1750
rect 860 -1765 910 -1750
rect 960 -1765 1010 -1750
rect 1060 -1765 1110 -1750
rect 335 -1920 395 -1910
rect 55 -1930 95 -1920
rect 55 -1945 65 -1930
rect 0 -1950 65 -1945
rect 85 -1945 95 -1930
rect 335 -1940 365 -1920
rect 385 -1930 755 -1920
rect 385 -1935 725 -1930
rect 385 -1940 395 -1935
rect 335 -1945 395 -1940
rect 85 -1950 150 -1945
rect 0 -1960 150 -1950
rect 0 -1975 50 -1960
rect 100 -1975 150 -1960
rect 200 -1950 395 -1945
rect 715 -1950 725 -1935
rect 745 -1945 755 -1930
rect 1015 -1930 1055 -1920
rect 1015 -1945 1025 -1930
rect 745 -1950 910 -1945
rect 200 -1960 350 -1950
rect 715 -1960 910 -1950
rect 200 -1975 250 -1960
rect 300 -1975 350 -1960
rect 480 -1975 530 -1960
rect 580 -1975 630 -1960
rect 760 -1975 810 -1960
rect 860 -1975 910 -1960
rect 960 -1950 1025 -1945
rect 1045 -1945 1055 -1930
rect 1045 -1950 1110 -1945
rect 960 -1960 1110 -1950
rect 960 -1975 1010 -1960
rect 1060 -1975 1110 -1960
rect 0 -2590 50 -2575
rect 100 -2590 150 -2575
rect 200 -2590 250 -2575
rect 300 -2590 350 -2575
rect 480 -2590 530 -2575
rect 580 -2590 630 -2575
rect 760 -2590 810 -2575
rect 860 -2590 910 -2575
rect 960 -2590 1010 -2575
rect 1060 -2590 1110 -2575
rect 480 -2600 630 -2590
rect 480 -2610 545 -2600
rect 535 -2620 545 -2610
rect 565 -2610 630 -2600
rect 565 -2620 575 -2610
rect 535 -2630 575 -2620
<< polycont >>
rect 880 640 900 660
rect -40 -30 -20 -10
rect 1130 -35 1150 -15
rect -40 -95 -20 -75
rect 65 -290 85 -270
rect 365 -290 385 -270
rect 545 -290 565 -270
rect 725 -290 745 -270
rect 1025 -290 1045 -270
rect 595 -1000 615 -980
rect 215 -1065 235 -1045
rect 485 -1065 505 -1045
rect 605 -1065 625 -1045
rect 1025 -1060 1045 -1040
rect 65 -1125 85 -1105
rect 365 -1125 385 -1105
rect 725 -1125 745 -1105
rect 1025 -1125 1045 -1105
rect 65 -1950 85 -1930
rect 365 -1940 385 -1920
rect 725 -1950 745 -1930
rect 1025 -1950 1045 -1930
rect 545 -2620 565 -2600
<< locali >>
rect 860 660 1210 670
rect 860 640 880 660
rect 900 640 1210 660
rect 860 630 1210 640
rect -95 600 -5 610
rect -95 30 -85 600
rect -65 30 -35 600
rect -15 30 -5 600
rect -95 20 -5 30
rect -50 -10 -5 20
rect -50 -30 -40 -10
rect -20 -30 -5 -10
rect -50 -40 -5 -30
rect 55 600 95 610
rect 55 30 65 600
rect 85 30 95 600
rect 55 -65 95 30
rect 155 600 195 610
rect 155 30 165 600
rect 185 30 195 600
rect 155 20 195 30
rect 255 600 295 610
rect 255 30 265 600
rect 285 30 295 600
rect -100 -75 95 -65
rect -100 -95 -40 -75
rect -20 -85 95 -75
rect -20 -95 -10 -85
rect -100 -105 -10 -95
rect 255 -125 295 30
rect 335 600 375 610
rect 335 30 345 600
rect 365 30 375 600
rect 335 -95 375 30
rect 435 600 475 610
rect 435 30 445 600
rect 465 30 475 600
rect 435 25 475 30
rect 535 600 575 610
rect 535 30 545 600
rect 565 30 575 600
rect 535 -45 575 30
rect 635 600 675 610
rect 635 30 645 600
rect 665 30 675 600
rect 635 25 675 30
rect 735 600 775 610
rect 735 30 745 600
rect 765 30 775 600
rect 535 -65 545 -45
rect 565 -65 575 -45
rect 535 -75 575 -65
rect 735 -85 775 30
rect 735 -95 745 -85
rect 335 -105 745 -95
rect 765 -105 775 -85
rect 335 -115 775 -105
rect 815 600 855 610
rect 815 30 825 600
rect 845 30 855 600
rect 255 -145 265 -125
rect 285 -135 295 -125
rect 815 -135 855 30
rect 915 600 955 610
rect 915 30 925 600
rect 945 30 955 600
rect 915 20 955 30
rect 1015 600 1055 630
rect 1015 30 1025 600
rect 1045 30 1055 600
rect 1015 20 1055 30
rect 1115 600 1205 610
rect 1115 30 1125 600
rect 1145 30 1175 600
rect 1195 30 1205 600
rect 1115 20 1205 30
rect 1115 -15 1160 20
rect 1115 -35 1130 -15
rect 1150 -35 1160 -15
rect 1115 -45 1160 -35
rect 285 -145 855 -135
rect 255 -155 855 -145
rect 355 -240 755 -220
rect -50 -270 95 -260
rect -50 -280 65 -270
rect -50 -320 -5 -280
rect -95 -330 -5 -320
rect -95 -900 -85 -330
rect -65 -900 -35 -330
rect -15 -900 -5 -330
rect -95 -910 -5 -900
rect 55 -290 65 -280
rect 85 -290 95 -270
rect 55 -330 95 -290
rect 355 -270 395 -240
rect 355 -290 365 -270
rect 385 -290 395 -270
rect 55 -900 65 -330
rect 85 -900 95 -330
rect 55 -910 95 -900
rect 155 -330 195 -320
rect 155 -900 165 -330
rect 185 -900 195 -330
rect 155 -910 195 -900
rect 255 -330 295 -320
rect 255 -900 265 -330
rect 285 -900 295 -330
rect 255 -930 295 -900
rect 355 -330 395 -290
rect 535 -270 575 -260
rect 535 -290 545 -270
rect 565 -290 575 -270
rect 355 -900 365 -330
rect 385 -900 395 -330
rect 355 -910 395 -900
rect 435 -330 475 -320
rect 435 -900 445 -330
rect 465 -900 475 -330
rect 435 -930 475 -900
rect 535 -330 575 -290
rect 715 -270 755 -240
rect 715 -290 725 -270
rect 745 -290 755 -270
rect 535 -900 545 -330
rect 565 -900 575 -330
rect 535 -910 575 -900
rect 635 -330 675 -320
rect 635 -900 645 -330
rect 665 -900 675 -330
rect 635 -930 675 -900
rect 715 -330 755 -290
rect 1015 -270 1160 -260
rect 1015 -290 1025 -270
rect 1045 -280 1160 -270
rect 1045 -290 1055 -280
rect 715 -900 725 -330
rect 745 -900 755 -330
rect 715 -910 755 -900
rect 815 -330 855 -320
rect 815 -900 825 -330
rect 845 -900 855 -330
rect 815 -930 855 -900
rect 915 -330 955 -320
rect 915 -900 925 -330
rect 945 -900 955 -330
rect 915 -910 955 -900
rect 1015 -330 1055 -290
rect 1015 -900 1025 -330
rect 1045 -900 1055 -330
rect 1015 -910 1055 -900
rect 1115 -320 1160 -280
rect 1115 -330 1205 -320
rect 1115 -900 1125 -330
rect 1145 -900 1175 -330
rect 1195 -900 1205 -330
rect 1115 -910 1205 -900
rect 255 -950 855 -930
rect 535 -980 1210 -970
rect 535 -1000 595 -980
rect 615 -990 1210 -980
rect 615 -1000 630 -990
rect 535 -1010 630 -1000
rect 200 -1045 250 -1035
rect 200 -1055 215 -1045
rect 155 -1065 215 -1055
rect 235 -1055 250 -1045
rect 475 -1045 515 -1035
rect 475 -1055 485 -1045
rect 235 -1065 485 -1055
rect 505 -1065 515 -1045
rect 155 -1075 515 -1065
rect -50 -1105 95 -1095
rect -50 -1115 65 -1105
rect -50 -1155 -5 -1115
rect -95 -1165 -5 -1155
rect -95 -1735 -85 -1165
rect -65 -1735 -35 -1165
rect -15 -1735 -5 -1165
rect -95 -1745 -5 -1735
rect 55 -1125 65 -1115
rect 85 -1125 95 -1105
rect 55 -1165 95 -1125
rect 55 -1735 65 -1165
rect 85 -1735 95 -1165
rect 55 -1745 95 -1735
rect 155 -1165 195 -1075
rect 355 -1105 395 -1095
rect 355 -1125 365 -1105
rect 385 -1125 395 -1105
rect 155 -1735 165 -1165
rect 185 -1735 195 -1165
rect 155 -1745 195 -1735
rect 255 -1165 295 -1155
rect 255 -1735 265 -1165
rect 285 -1735 295 -1165
rect 255 -1765 295 -1735
rect 355 -1165 395 -1125
rect 355 -1735 365 -1165
rect 385 -1735 395 -1165
rect 355 -1745 395 -1735
rect 435 -1165 475 -1155
rect 435 -1735 445 -1165
rect 465 -1735 475 -1165
rect 435 -1765 475 -1735
rect 535 -1165 575 -1010
rect 595 -1045 635 -1035
rect 595 -1065 605 -1045
rect 625 -1055 635 -1045
rect 1015 -1040 1055 -1030
rect 625 -1065 955 -1055
rect 595 -1075 955 -1065
rect 1015 -1060 1025 -1040
rect 1045 -1050 1055 -1040
rect 1045 -1060 1210 -1050
rect 1015 -1070 1210 -1060
rect 715 -1105 755 -1095
rect 715 -1125 725 -1105
rect 745 -1125 755 -1105
rect 535 -1735 545 -1165
rect 565 -1735 575 -1165
rect 535 -1745 575 -1735
rect 635 -1165 675 -1155
rect 635 -1735 645 -1165
rect 665 -1735 675 -1165
rect 635 -1765 675 -1735
rect 715 -1165 755 -1125
rect 715 -1735 725 -1165
rect 745 -1735 755 -1165
rect 715 -1745 755 -1735
rect 815 -1165 855 -1155
rect 815 -1735 825 -1165
rect 845 -1735 855 -1165
rect 815 -1765 855 -1735
rect 915 -1165 955 -1075
rect 915 -1735 925 -1165
rect 945 -1735 955 -1165
rect 915 -1745 955 -1735
rect 1015 -1105 1160 -1095
rect 1015 -1125 1025 -1105
rect 1045 -1115 1160 -1105
rect 1045 -1125 1055 -1115
rect 1015 -1165 1055 -1125
rect 1015 -1735 1025 -1165
rect 1045 -1735 1055 -1165
rect 1015 -1745 1055 -1735
rect 1115 -1155 1160 -1115
rect 1115 -1165 1205 -1155
rect 1115 -1735 1125 -1165
rect 1145 -1735 1175 -1165
rect 1195 -1735 1205 -1165
rect 1115 -1745 1205 -1735
rect 255 -1805 855 -1765
rect 255 -1845 855 -1825
rect -50 -1930 95 -1920
rect -50 -1940 65 -1930
rect -50 -1980 -5 -1940
rect 55 -1950 65 -1940
rect 85 -1950 95 -1930
rect 55 -1960 95 -1950
rect -95 -1990 -5 -1980
rect -95 -2560 -85 -1990
rect -65 -2560 -35 -1990
rect -15 -2560 -5 -1990
rect -95 -2570 -5 -2560
rect 55 -1990 95 -1980
rect 55 -2560 65 -1990
rect 85 -2560 95 -1990
rect 55 -2570 95 -2560
rect 155 -1990 195 -1980
rect 155 -2560 165 -1990
rect 185 -2560 195 -1990
rect 155 -2570 195 -2560
rect 255 -1990 295 -1845
rect 255 -2560 265 -1990
rect 285 -2560 295 -1990
rect 255 -2570 295 -2560
rect 355 -1920 395 -1910
rect 355 -1940 365 -1920
rect 385 -1940 395 -1920
rect 355 -1990 395 -1940
rect 355 -2560 365 -1990
rect 385 -2560 395 -1990
rect 355 -2570 395 -2560
rect 435 -1990 475 -1845
rect 435 -2560 445 -1990
rect 465 -2560 475 -1990
rect 435 -2570 475 -2560
rect 535 -1875 575 -1865
rect 535 -1895 545 -1875
rect 565 -1895 575 -1875
rect 535 -1990 575 -1895
rect 535 -2560 545 -1990
rect 565 -2560 575 -1990
rect 535 -2600 575 -2560
rect 635 -1990 675 -1845
rect 635 -2560 645 -1990
rect 665 -2560 675 -1990
rect 635 -2570 675 -2560
rect 715 -1930 755 -1920
rect 715 -1950 725 -1930
rect 745 -1950 755 -1930
rect 715 -1990 755 -1950
rect 715 -2560 725 -1990
rect 745 -2560 755 -1990
rect 715 -2570 755 -2560
rect 815 -1990 855 -1845
rect 1015 -1930 1160 -1920
rect 1015 -1950 1025 -1930
rect 1045 -1945 1160 -1930
rect 1045 -1950 1055 -1945
rect 815 -2560 825 -1990
rect 845 -2560 855 -1990
rect 815 -2570 855 -2560
rect 915 -1990 955 -1980
rect 915 -2560 925 -1990
rect 945 -2560 955 -1990
rect 915 -2570 955 -2560
rect 1015 -1990 1055 -1950
rect 1015 -2560 1025 -1990
rect 1045 -2560 1055 -1990
rect 1015 -2570 1055 -2560
rect 1115 -1980 1160 -1945
rect 1115 -1990 1205 -1980
rect 1115 -2560 1125 -1990
rect 1145 -2560 1175 -1990
rect 1195 -2560 1205 -1990
rect 1115 -2570 1205 -2560
rect 535 -2620 545 -2600
rect 565 -2610 575 -2600
rect 565 -2620 1210 -2610
rect 535 -2630 1210 -2620
<< viali >>
rect -85 30 -65 600
rect -35 30 -15 600
rect 165 30 185 600
rect 445 30 465 600
rect 645 30 665 600
rect 545 -65 565 -45
rect 745 -105 765 -85
rect 265 -145 285 -125
rect 925 30 945 600
rect 1125 30 1145 600
rect 1175 30 1195 600
rect -85 -900 -65 -330
rect -35 -900 -15 -330
rect 65 -900 85 -330
rect 165 -900 185 -330
rect 925 -900 945 -330
rect 1025 -900 1045 -330
rect 1125 -900 1145 -330
rect 1175 -900 1195 -330
rect -85 -1735 -65 -1165
rect -35 -1735 -15 -1165
rect 65 -1735 85 -1165
rect 365 -1125 385 -1105
rect 265 -1735 285 -1165
rect 825 -1735 845 -1165
rect 1025 -1735 1045 -1165
rect 1125 -1735 1145 -1165
rect 1175 -1735 1195 -1165
rect -85 -2560 -65 -1990
rect -35 -2560 -15 -1990
rect 65 -2560 85 -1990
rect 165 -2560 185 -1990
rect 365 -1940 385 -1920
rect 545 -1895 565 -1875
rect 925 -2560 945 -1990
rect 1025 -2560 1045 -1990
rect 1125 -2560 1145 -1990
rect 1175 -2560 1195 -1990
<< metal1 >>
rect -100 600 1210 610
rect -100 30 -85 600
rect -65 30 -35 600
rect -15 30 165 600
rect 185 30 445 600
rect 465 30 645 600
rect 665 30 925 600
rect 945 30 1125 600
rect 1145 30 1175 600
rect 1195 30 1210 600
rect -100 20 1210 30
rect -100 -330 195 20
rect 535 -45 575 -35
rect 535 -65 545 -45
rect 565 -65 575 -45
rect -100 -900 -85 -330
rect -65 -900 -35 -330
rect -15 -900 65 -330
rect 85 -900 165 -330
rect 185 -900 195 -330
rect -100 -910 195 -900
rect 255 -125 295 -115
rect 255 -145 265 -125
rect 285 -145 295 -125
rect 255 -1095 295 -145
rect 255 -1105 395 -1095
rect 255 -1125 365 -1105
rect 385 -1125 395 -1105
rect 355 -1135 395 -1125
rect -100 -1165 300 -1155
rect -100 -1735 -85 -1165
rect -65 -1735 -35 -1165
rect -15 -1735 65 -1165
rect 85 -1735 265 -1165
rect 285 -1735 300 -1165
rect -100 -1980 300 -1735
rect 535 -1765 575 -65
rect 355 -1805 575 -1765
rect 735 -85 775 -75
rect 735 -105 745 -85
rect 765 -105 775 -85
rect 355 -1920 395 -1805
rect 735 -1865 775 -105
rect 915 -330 1210 20
rect 915 -900 925 -330
rect 945 -900 1025 -330
rect 1045 -900 1125 -330
rect 1145 -900 1175 -330
rect 1195 -900 1210 -330
rect 915 -910 1210 -900
rect 535 -1875 775 -1865
rect 535 -1895 545 -1875
rect 565 -1895 775 -1875
rect 535 -1905 775 -1895
rect 810 -1165 1210 -1155
rect 810 -1735 825 -1165
rect 845 -1735 1025 -1165
rect 1045 -1735 1125 -1165
rect 1145 -1735 1175 -1165
rect 1195 -1735 1210 -1165
rect 355 -1940 365 -1920
rect 385 -1940 395 -1920
rect 355 -1950 395 -1940
rect 810 -1980 1210 -1735
rect -100 -1990 1210 -1980
rect -100 -2560 -85 -1990
rect -65 -2560 -35 -1990
rect -15 -2560 65 -1990
rect 85 -2560 165 -1990
rect 185 -2560 925 -1990
rect 945 -2560 1025 -1990
rect 1045 -2560 1125 -1990
rect 1145 -2560 1175 -1990
rect 1195 -2560 1210 -1990
rect -100 -2570 1210 -2560
<< labels >>
rlabel locali 1210 -2620 1210 -2620 3 Vcn
rlabel metal1 -100 -2275 -100 -2275 7 VN
rlabel locali 1210 -980 1210 -980 3 Vcp
rlabel metal1 -100 315 -100 315 7 VP
rlabel locali -100 -85 -100 -85 7 Vbp
rlabel locali 1210 -1060 1210 -1060 3 Vbn
<< end >>
