magic
tech sky130A
timestamp 1615581013
<< nmos >>
rect -15 620 35 770
rect 85 620 135 770
rect 185 620 235 770
rect 285 620 335 770
rect 385 620 435 770
rect 485 620 535 770
rect 585 620 635 770
rect 685 620 735 770
rect 785 620 835 770
rect 885 620 935 770
rect -15 79 35 379
rect 85 79 135 379
rect 185 79 235 379
rect 285 79 335 379
rect 385 79 435 379
rect 485 79 535 379
rect 585 79 635 379
rect 685 79 735 379
rect 785 79 835 379
rect 885 79 935 379
rect -15 -765 35 -165
rect 85 -765 135 -165
rect 185 -765 235 -165
rect 285 -765 335 -165
rect 385 -765 435 -165
rect 485 -765 535 -165
rect 585 -765 635 -165
rect 685 -765 735 -165
rect 785 -765 835 -165
rect 885 -765 935 -165
rect -15 -1665 35 -1065
rect 85 -1665 135 -1065
rect 185 -1665 235 -1065
rect 285 -1665 335 -1065
rect 385 -1665 435 -1065
rect 485 -1665 535 -1065
rect 585 -1665 635 -1065
rect 685 -1665 735 -1065
rect 785 -1665 835 -1065
rect 885 -1665 935 -1065
<< ndiff >>
rect -65 760 -15 770
rect -65 635 -50 760
rect -30 635 -15 760
rect -65 620 -15 635
rect 35 760 85 770
rect 35 635 50 760
rect 70 635 85 760
rect 35 620 85 635
rect 135 760 185 770
rect 135 635 150 760
rect 170 635 185 760
rect 135 620 185 635
rect 235 760 285 770
rect 235 635 250 760
rect 270 635 285 760
rect 235 620 285 635
rect 335 760 385 770
rect 335 635 350 760
rect 370 635 385 760
rect 335 620 385 635
rect 435 760 485 770
rect 435 635 450 760
rect 470 635 485 760
rect 435 620 485 635
rect 535 760 585 770
rect 535 635 550 760
rect 570 635 585 760
rect 535 620 585 635
rect 635 760 685 770
rect 635 635 650 760
rect 670 635 685 760
rect 635 620 685 635
rect 735 760 785 770
rect 735 635 750 760
rect 770 635 785 760
rect 735 620 785 635
rect 835 760 885 770
rect 835 635 850 760
rect 870 635 885 760
rect 835 620 885 635
rect 935 760 985 770
rect 935 635 950 760
rect 970 635 985 760
rect 935 620 985 635
rect -65 364 -15 379
rect -65 94 -50 364
rect -30 94 -15 364
rect -65 79 -15 94
rect 35 364 85 379
rect 35 94 50 364
rect 70 94 85 364
rect 35 79 85 94
rect 135 364 185 379
rect 135 94 150 364
rect 170 94 185 364
rect 135 79 185 94
rect 235 364 285 379
rect 235 94 250 364
rect 270 94 285 364
rect 235 79 285 94
rect 335 364 385 379
rect 335 94 350 364
rect 370 94 385 364
rect 335 79 385 94
rect 435 364 485 379
rect 435 94 450 364
rect 470 94 485 364
rect 435 79 485 94
rect 535 364 585 379
rect 535 94 550 364
rect 570 94 585 364
rect 535 79 585 94
rect 635 364 685 379
rect 635 94 650 364
rect 670 94 685 364
rect 635 79 685 94
rect 735 364 785 379
rect 735 94 750 364
rect 770 94 785 364
rect 735 79 785 94
rect 835 364 885 379
rect 835 94 850 364
rect 870 94 885 364
rect 835 79 885 94
rect 935 364 985 379
rect 935 94 950 364
rect 970 94 985 364
rect 935 79 985 94
rect -65 -180 -15 -165
rect -65 -750 -50 -180
rect -30 -750 -15 -180
rect -65 -765 -15 -750
rect 35 -180 85 -165
rect 35 -750 50 -180
rect 70 -750 85 -180
rect 35 -765 85 -750
rect 135 -180 185 -165
rect 135 -750 150 -180
rect 170 -750 185 -180
rect 135 -765 185 -750
rect 235 -180 285 -165
rect 235 -750 250 -180
rect 270 -750 285 -180
rect 235 -765 285 -750
rect 335 -180 385 -165
rect 335 -750 350 -180
rect 370 -750 385 -180
rect 335 -765 385 -750
rect 435 -180 485 -165
rect 435 -750 450 -180
rect 470 -750 485 -180
rect 435 -765 485 -750
rect 535 -180 585 -165
rect 535 -750 550 -180
rect 570 -750 585 -180
rect 535 -765 585 -750
rect 635 -180 685 -165
rect 635 -750 650 -180
rect 670 -750 685 -180
rect 635 -765 685 -750
rect 735 -180 785 -165
rect 735 -750 750 -180
rect 770 -750 785 -180
rect 735 -765 785 -750
rect 835 -180 885 -165
rect 835 -750 850 -180
rect 870 -750 885 -180
rect 835 -765 885 -750
rect 935 -180 985 -165
rect 935 -750 950 -180
rect 970 -750 985 -180
rect 935 -765 985 -750
rect -65 -1080 -15 -1065
rect -65 -1650 -50 -1080
rect -30 -1650 -15 -1080
rect -65 -1665 -15 -1650
rect 35 -1080 85 -1065
rect 35 -1650 50 -1080
rect 70 -1650 85 -1080
rect 35 -1665 85 -1650
rect 135 -1080 185 -1065
rect 135 -1650 150 -1080
rect 170 -1650 185 -1080
rect 135 -1665 185 -1650
rect 235 -1080 285 -1065
rect 235 -1650 250 -1080
rect 270 -1650 285 -1080
rect 235 -1665 285 -1650
rect 335 -1080 385 -1065
rect 335 -1650 350 -1080
rect 370 -1650 385 -1080
rect 335 -1665 385 -1650
rect 435 -1080 485 -1065
rect 435 -1650 450 -1080
rect 470 -1650 485 -1080
rect 435 -1665 485 -1650
rect 535 -1080 585 -1065
rect 535 -1650 550 -1080
rect 570 -1650 585 -1080
rect 535 -1665 585 -1650
rect 635 -1080 685 -1065
rect 635 -1650 650 -1080
rect 670 -1650 685 -1080
rect 635 -1665 685 -1650
rect 735 -1080 785 -1065
rect 735 -1650 750 -1080
rect 770 -1650 785 -1080
rect 735 -1665 785 -1650
rect 835 -1080 885 -1065
rect 835 -1650 850 -1080
rect 870 -1650 885 -1080
rect 835 -1665 885 -1650
rect 935 -1080 985 -1065
rect 935 -1650 950 -1080
rect 970 -1650 985 -1080
rect 935 -1665 985 -1650
<< ndiffc >>
rect -50 635 -30 760
rect 50 635 70 760
rect 150 635 170 760
rect 250 635 270 760
rect 350 635 370 760
rect 450 635 470 760
rect 550 635 570 760
rect 650 635 670 760
rect 750 635 770 760
rect 850 635 870 760
rect 950 635 970 760
rect -50 94 -30 364
rect 50 94 70 364
rect 150 94 170 364
rect 250 94 270 364
rect 350 94 370 364
rect 450 94 470 364
rect 550 94 570 364
rect 650 94 670 364
rect 750 94 770 364
rect 850 94 870 364
rect 950 94 970 364
rect -50 -750 -30 -180
rect 50 -750 70 -180
rect 150 -750 170 -180
rect 250 -750 270 -180
rect 350 -750 370 -180
rect 450 -750 470 -180
rect 550 -750 570 -180
rect 650 -750 670 -180
rect 750 -750 770 -180
rect 850 -750 870 -180
rect 950 -750 970 -180
rect -50 -1650 -30 -1080
rect 50 -1650 70 -1080
rect 150 -1650 170 -1080
rect 250 -1650 270 -1080
rect 350 -1650 370 -1080
rect 450 -1650 470 -1080
rect 550 -1650 570 -1080
rect 650 -1650 670 -1080
rect 750 -1650 770 -1080
rect 850 -1650 870 -1080
rect 950 -1650 970 -1080
<< psubdiff >>
rect -115 760 -65 770
rect -115 635 -100 760
rect -80 635 -65 760
rect -115 620 -65 635
rect 985 760 1035 770
rect 985 635 1000 760
rect 1020 635 1035 760
rect 985 620 1035 635
rect -115 364 -65 379
rect -115 94 -100 364
rect -80 94 -65 364
rect -115 79 -65 94
rect 985 364 1035 379
rect 985 94 1000 364
rect 1020 94 1035 364
rect 985 79 1035 94
rect -115 -180 -65 -165
rect -115 -750 -100 -180
rect -80 -750 -65 -180
rect -115 -765 -65 -750
rect 985 -180 1035 -165
rect 985 -750 1000 -180
rect 1020 -750 1035 -180
rect 985 -765 1035 -750
rect -115 -1080 -65 -1065
rect -115 -1650 -100 -1080
rect -80 -1650 -65 -1080
rect -115 -1665 -65 -1650
rect 985 -1080 1035 -1065
rect 985 -1650 1000 -1080
rect 1020 -1650 1035 -1080
rect 985 -1665 1035 -1650
<< psubdiffcont >>
rect -100 635 -80 760
rect 1000 635 1020 760
rect -100 94 -80 364
rect 1000 94 1020 364
rect -100 -750 -80 -180
rect 1000 -750 1020 -180
rect -100 -1650 -80 -1080
rect 1000 -1650 1020 -1080
<< poly >>
rect -15 770 35 785
rect 85 770 135 785
rect 185 770 235 785
rect 285 770 335 785
rect 385 770 435 785
rect 485 770 535 785
rect 585 770 635 785
rect 685 770 735 785
rect 785 770 835 785
rect 885 770 935 785
rect -15 610 35 620
rect 85 610 135 620
rect 185 610 235 620
rect 285 610 335 620
rect 385 610 435 620
rect 485 610 535 620
rect 585 610 635 620
rect 685 610 735 620
rect 785 610 835 620
rect -60 600 35 610
rect -60 580 -50 600
rect -30 595 35 600
rect 60 595 835 610
rect 885 610 935 620
rect 885 600 980 610
rect 885 595 950 600
rect -30 580 -20 595
rect -60 570 -20 580
rect 60 545 75 595
rect 940 580 950 595
rect 970 580 980 600
rect 940 570 980 580
rect -65 535 75 545
rect -65 515 -55 535
rect -35 530 75 535
rect -35 515 -25 530
rect -65 505 -25 515
rect -15 379 35 394
rect 85 379 135 394
rect 185 379 235 394
rect 285 379 335 394
rect 385 379 435 394
rect 485 379 535 394
rect 585 379 635 394
rect 685 379 735 394
rect 785 379 835 394
rect 885 379 935 394
rect -15 64 35 79
rect 85 64 135 79
rect 185 64 235 79
rect 285 64 335 79
rect 385 64 435 79
rect 485 64 535 79
rect 585 64 635 79
rect 685 64 735 79
rect 785 64 835 79
rect 885 64 935 79
rect -15 -165 35 -150
rect 85 -165 135 -150
rect 185 -165 235 -150
rect 285 -165 335 -150
rect 385 -165 435 -150
rect 485 -165 535 -150
rect 585 -165 635 -150
rect 685 -165 735 -150
rect 785 -165 835 -150
rect 885 -165 935 -150
rect -15 -780 35 -765
rect 85 -780 135 -765
rect 185 -780 235 -765
rect 285 -780 335 -765
rect 385 -780 435 -765
rect 485 -780 535 -765
rect 585 -780 635 -765
rect 685 -780 735 -765
rect 785 -780 835 -765
rect 885 -780 935 -765
rect -15 -1065 35 -1050
rect 85 -1065 135 -1050
rect 185 -1065 235 -1050
rect 285 -1065 335 -1050
rect 385 -1065 435 -1050
rect 485 -1065 535 -1050
rect 585 -1065 635 -1050
rect 685 -1065 735 -1050
rect 785 -1065 835 -1050
rect 885 -1065 935 -1050
rect -15 -1680 35 -1665
rect 85 -1680 135 -1665
rect 185 -1680 235 -1665
rect 285 -1680 335 -1665
rect 385 -1680 435 -1665
rect 485 -1680 535 -1665
rect 585 -1680 635 -1665
rect 685 -1680 735 -1665
rect 785 -1680 835 -1665
rect 885 -1680 935 -1665
<< polycont >>
rect -50 580 -30 600
rect 950 580 970 600
rect -55 515 -35 535
<< locali >>
rect -110 760 -20 765
rect -110 635 -100 760
rect -80 635 -50 760
rect -30 635 -20 760
rect -110 625 -20 635
rect 40 760 80 765
rect 40 635 50 760
rect 70 635 80 760
rect 40 625 80 635
rect 140 760 180 765
rect 140 635 150 760
rect 170 635 180 760
rect 140 625 180 635
rect 240 760 280 765
rect 240 635 250 760
rect 270 635 280 760
rect 240 625 280 635
rect 340 760 380 765
rect 340 635 350 760
rect 370 635 380 760
rect 340 625 380 635
rect 440 760 480 765
rect 440 635 450 760
rect 470 635 480 760
rect 440 625 480 635
rect 540 760 580 765
rect 540 635 550 760
rect 570 635 580 760
rect 540 625 580 635
rect 640 760 680 765
rect 640 635 650 760
rect 670 635 680 760
rect 640 625 680 635
rect 740 760 780 765
rect 740 635 750 760
rect 770 635 780 760
rect 740 625 780 635
rect 840 760 880 765
rect 840 635 850 760
rect 870 635 880 760
rect 840 625 880 635
rect 940 760 1030 765
rect 940 635 950 760
rect 970 635 1000 760
rect 1020 635 1030 760
rect 940 625 1030 635
rect -60 600 -20 625
rect -60 580 -50 600
rect -30 580 -20 600
rect -60 570 -20 580
rect 940 600 980 625
rect 940 580 950 600
rect 970 580 980 600
rect 940 570 980 580
rect -115 535 -25 545
rect -115 525 -55 535
rect -65 515 -55 525
rect -35 515 -25 535
rect -65 505 -25 515
rect -110 364 -20 374
rect -110 94 -100 364
rect -80 94 -50 364
rect -30 94 -20 364
rect -110 84 -20 94
rect 40 364 80 374
rect 40 94 50 364
rect 70 94 80 364
rect 40 84 80 94
rect 140 364 180 374
rect 140 94 150 364
rect 170 94 180 364
rect 140 84 180 94
rect 240 364 280 374
rect 240 94 250 364
rect 270 94 280 364
rect 240 84 280 94
rect 340 364 380 374
rect 340 94 350 364
rect 370 94 380 364
rect 340 84 380 94
rect 440 364 480 374
rect 440 94 450 364
rect 470 94 480 364
rect 440 84 480 94
rect 540 364 580 374
rect 540 94 550 364
rect 570 94 580 364
rect 540 84 580 94
rect 640 364 680 374
rect 640 94 650 364
rect 670 94 680 364
rect 640 84 680 94
rect 740 364 780 374
rect 740 94 750 364
rect 770 94 780 364
rect 740 84 780 94
rect 840 364 880 374
rect 840 94 850 364
rect 870 94 880 364
rect 840 84 880 94
rect 940 364 1030 374
rect 940 94 950 364
rect 970 94 1000 364
rect 1020 94 1030 364
rect 940 84 1030 94
rect -110 -180 -20 -170
rect -110 -750 -100 -180
rect -80 -750 -50 -180
rect -30 -750 -20 -180
rect -110 -760 -20 -750
rect 40 -180 80 -170
rect 40 -750 50 -180
rect 70 -750 80 -180
rect 40 -760 80 -750
rect 140 -180 180 -170
rect 140 -750 150 -180
rect 170 -750 180 -180
rect 140 -760 180 -750
rect 240 -180 280 -170
rect 240 -750 250 -180
rect 270 -750 280 -180
rect 240 -760 280 -750
rect 340 -180 380 -170
rect 340 -750 350 -180
rect 370 -750 380 -180
rect 340 -760 380 -750
rect 440 -180 480 -170
rect 440 -750 450 -180
rect 470 -750 480 -180
rect 440 -760 480 -750
rect 540 -180 580 -170
rect 540 -750 550 -180
rect 570 -750 580 -180
rect 540 -760 580 -750
rect 640 -180 680 -170
rect 640 -750 650 -180
rect 670 -750 680 -180
rect 640 -760 680 -750
rect 740 -180 780 -170
rect 740 -750 750 -180
rect 770 -750 780 -180
rect 740 -760 780 -750
rect 840 -180 880 -170
rect 840 -750 850 -180
rect 870 -750 880 -180
rect 840 -760 880 -750
rect 940 -180 1030 -170
rect 940 -750 950 -180
rect 970 -750 1000 -180
rect 1020 -750 1030 -180
rect 940 -760 1030 -750
rect -110 -1080 -20 -1070
rect -110 -1650 -100 -1080
rect -80 -1650 -50 -1080
rect -30 -1650 -20 -1080
rect -110 -1660 -20 -1650
rect 40 -1080 80 -1070
rect 40 -1650 50 -1080
rect 70 -1650 80 -1080
rect 40 -1660 80 -1650
rect 140 -1080 180 -1070
rect 140 -1650 150 -1080
rect 170 -1650 180 -1080
rect 140 -1660 180 -1650
rect 240 -1080 280 -1070
rect 240 -1650 250 -1080
rect 270 -1650 280 -1080
rect 240 -1660 280 -1650
rect 340 -1080 380 -1070
rect 340 -1650 350 -1080
rect 370 -1650 380 -1080
rect 340 -1660 380 -1650
rect 440 -1080 480 -1070
rect 440 -1650 450 -1080
rect 470 -1650 480 -1080
rect 440 -1660 480 -1650
rect 540 -1080 580 -1070
rect 540 -1650 550 -1080
rect 570 -1650 580 -1080
rect 540 -1660 580 -1650
rect 640 -1080 680 -1070
rect 640 -1650 650 -1080
rect 670 -1650 680 -1080
rect 640 -1660 680 -1650
rect 740 -1080 780 -1070
rect 740 -1650 750 -1080
rect 770 -1650 780 -1080
rect 740 -1660 780 -1650
rect 840 -1080 880 -1070
rect 840 -1650 850 -1080
rect 870 -1650 880 -1080
rect 840 -1660 880 -1650
rect 940 -1080 1030 -1070
rect 940 -1650 950 -1080
rect 970 -1650 1000 -1080
rect 1020 -1650 1030 -1080
rect 940 -1660 1030 -1650
<< end >>
