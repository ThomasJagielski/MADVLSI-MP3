magic
tech sky130A
timestamp 1615643413
<< nwell >>
rect -135 -830 1055 795
<< nmos >>
rect -15 -1765 35 -1165
rect 85 -1765 135 -1165
rect 185 -1765 235 -1165
rect 285 -1765 335 -1165
rect 385 -1765 435 -1165
rect 485 -1765 535 -1165
rect 585 -1765 635 -1165
rect 685 -1765 735 -1165
rect 785 -1765 835 -1165
rect 885 -1765 935 -1165
<< pmos >>
rect -15 625 35 775
rect 85 625 135 775
rect 185 625 235 775
rect 285 625 335 775
rect 385 625 435 775
rect 485 625 535 775
rect 585 625 635 775
rect 685 625 735 775
rect 785 625 835 775
rect 885 625 935 775
rect -15 80 35 380
rect 85 80 135 380
rect 185 80 235 380
rect 285 80 335 380
rect 385 80 435 380
rect 485 80 535 380
rect 585 80 635 380
rect 685 80 735 380
rect 785 80 835 380
rect 885 80 935 380
rect -15 -810 35 -210
rect 85 -810 135 -210
rect 185 -810 235 -210
rect 285 -810 335 -210
rect 385 -810 435 -210
rect 485 -810 535 -210
rect 585 -810 635 -210
rect 685 -810 735 -210
rect 785 -810 835 -210
rect 885 -810 935 -210
<< ndiff >>
rect -65 -1180 -15 -1165
rect -65 -1750 -50 -1180
rect -30 -1750 -15 -1180
rect -65 -1765 -15 -1750
rect 35 -1180 85 -1165
rect 35 -1750 50 -1180
rect 70 -1750 85 -1180
rect 35 -1765 85 -1750
rect 135 -1180 185 -1165
rect 135 -1750 150 -1180
rect 170 -1750 185 -1180
rect 135 -1765 185 -1750
rect 235 -1180 285 -1165
rect 235 -1750 250 -1180
rect 270 -1750 285 -1180
rect 235 -1765 285 -1750
rect 335 -1180 385 -1165
rect 335 -1750 350 -1180
rect 370 -1750 385 -1180
rect 335 -1765 385 -1750
rect 435 -1180 485 -1165
rect 435 -1750 450 -1180
rect 470 -1750 485 -1180
rect 435 -1765 485 -1750
rect 535 -1180 585 -1165
rect 535 -1750 550 -1180
rect 570 -1750 585 -1180
rect 535 -1765 585 -1750
rect 635 -1180 685 -1165
rect 635 -1750 650 -1180
rect 670 -1750 685 -1180
rect 635 -1765 685 -1750
rect 735 -1180 785 -1165
rect 735 -1750 750 -1180
rect 770 -1750 785 -1180
rect 735 -1765 785 -1750
rect 835 -1180 885 -1165
rect 835 -1750 850 -1180
rect 870 -1750 885 -1180
rect 835 -1765 885 -1750
rect 935 -1180 985 -1165
rect 935 -1750 950 -1180
rect 970 -1750 985 -1180
rect 935 -1765 985 -1750
<< pdiff >>
rect -65 765 -15 775
rect -65 640 -50 765
rect -30 640 -15 765
rect -65 625 -15 640
rect 35 765 85 775
rect 35 640 50 765
rect 70 640 85 765
rect 35 625 85 640
rect 135 765 185 775
rect 135 640 150 765
rect 170 640 185 765
rect 135 625 185 640
rect 235 765 285 775
rect 235 640 250 765
rect 270 640 285 765
rect 235 625 285 640
rect 335 765 385 775
rect 335 640 350 765
rect 370 640 385 765
rect 335 625 385 640
rect 435 765 485 775
rect 435 640 450 765
rect 470 640 485 765
rect 435 625 485 640
rect 535 765 585 775
rect 535 640 550 765
rect 570 640 585 765
rect 535 625 585 640
rect 635 765 685 775
rect 635 640 650 765
rect 670 640 685 765
rect 635 625 685 640
rect 735 765 785 775
rect 735 640 750 765
rect 770 640 785 765
rect 735 625 785 640
rect 835 765 885 775
rect 835 640 850 765
rect 870 640 885 765
rect 835 625 885 640
rect 935 765 985 775
rect 935 640 950 765
rect 970 640 985 765
rect 935 625 985 640
rect -65 365 -15 380
rect -65 95 -50 365
rect -30 95 -15 365
rect -65 80 -15 95
rect 35 365 85 380
rect 35 95 50 365
rect 70 95 85 365
rect 35 80 85 95
rect 135 365 185 380
rect 135 95 150 365
rect 170 95 185 365
rect 135 80 185 95
rect 235 365 285 380
rect 235 95 250 365
rect 270 95 285 365
rect 235 80 285 95
rect 335 365 385 380
rect 335 95 350 365
rect 370 95 385 365
rect 335 80 385 95
rect 435 365 485 380
rect 435 95 450 365
rect 470 95 485 365
rect 435 80 485 95
rect 535 365 585 380
rect 535 95 550 365
rect 570 95 585 365
rect 535 80 585 95
rect 635 365 685 380
rect 635 95 650 365
rect 670 95 685 365
rect 635 80 685 95
rect 735 365 785 380
rect 735 95 750 365
rect 770 95 785 365
rect 735 80 785 95
rect 835 365 885 380
rect 835 95 850 365
rect 870 95 885 365
rect 835 80 885 95
rect 935 365 985 380
rect 935 95 950 365
rect 970 95 985 365
rect 935 80 985 95
rect -65 -225 -15 -210
rect -65 -795 -50 -225
rect -30 -795 -15 -225
rect -65 -810 -15 -795
rect 35 -225 85 -210
rect 35 -795 50 -225
rect 70 -795 85 -225
rect 35 -810 85 -795
rect 135 -225 185 -210
rect 135 -795 150 -225
rect 170 -795 185 -225
rect 135 -810 185 -795
rect 235 -225 285 -210
rect 235 -795 250 -225
rect 270 -795 285 -225
rect 235 -810 285 -795
rect 335 -225 385 -210
rect 335 -795 350 -225
rect 370 -795 385 -225
rect 335 -810 385 -795
rect 435 -225 485 -210
rect 435 -795 450 -225
rect 470 -795 485 -225
rect 435 -810 485 -795
rect 535 -225 585 -210
rect 535 -795 550 -225
rect 570 -795 585 -225
rect 535 -810 585 -795
rect 635 -225 685 -210
rect 635 -795 650 -225
rect 670 -795 685 -225
rect 635 -810 685 -795
rect 735 -225 785 -210
rect 735 -795 750 -225
rect 770 -795 785 -225
rect 735 -810 785 -795
rect 835 -225 885 -210
rect 835 -795 850 -225
rect 870 -795 885 -225
rect 835 -810 885 -795
rect 935 -225 985 -210
rect 935 -795 950 -225
rect 970 -795 985 -225
rect 935 -810 985 -795
<< ndiffc >>
rect -50 -1750 -30 -1180
rect 50 -1750 70 -1180
rect 150 -1750 170 -1180
rect 250 -1750 270 -1180
rect 350 -1750 370 -1180
rect 450 -1750 470 -1180
rect 550 -1750 570 -1180
rect 650 -1750 670 -1180
rect 750 -1750 770 -1180
rect 850 -1750 870 -1180
rect 950 -1750 970 -1180
<< pdiffc >>
rect -50 640 -30 765
rect 50 640 70 765
rect 150 640 170 765
rect 250 640 270 765
rect 350 640 370 765
rect 450 640 470 765
rect 550 640 570 765
rect 650 640 670 765
rect 750 640 770 765
rect 850 640 870 765
rect 950 640 970 765
rect -50 95 -30 365
rect 50 95 70 365
rect 150 95 170 365
rect 250 95 270 365
rect 350 95 370 365
rect 450 95 470 365
rect 550 95 570 365
rect 650 95 670 365
rect 750 95 770 365
rect 850 95 870 365
rect 950 95 970 365
rect -50 -795 -30 -225
rect 50 -795 70 -225
rect 150 -795 170 -225
rect 250 -795 270 -225
rect 350 -795 370 -225
rect 450 -795 470 -225
rect 550 -795 570 -225
rect 650 -795 670 -225
rect 750 -795 770 -225
rect 850 -795 870 -225
rect 950 -795 970 -225
<< psubdiff >>
rect -115 -1180 -65 -1165
rect -115 -1750 -100 -1180
rect -80 -1750 -65 -1180
rect -115 -1765 -65 -1750
rect 985 -1180 1035 -1165
rect 985 -1750 1000 -1180
rect 1020 -1750 1035 -1180
rect 985 -1765 1035 -1750
<< nsubdiff >>
rect -115 765 -65 775
rect -115 640 -100 765
rect -80 640 -65 765
rect -115 625 -65 640
rect 985 765 1035 775
rect 985 640 1000 765
rect 1020 640 1035 765
rect 985 625 1035 640
rect -115 365 -65 380
rect -115 95 -100 365
rect -80 95 -65 365
rect -115 80 -65 95
rect 985 365 1035 380
rect 985 95 1000 365
rect 1020 95 1035 365
rect 985 80 1035 95
rect -115 -225 -65 -210
rect -115 -795 -100 -225
rect -80 -795 -65 -225
rect -115 -810 -65 -795
rect 985 -225 1035 -210
rect 985 -795 1000 -225
rect 1020 -795 1035 -225
rect 985 -810 1035 -795
<< psubdiffcont >>
rect -100 -1750 -80 -1180
rect 1000 -1750 1020 -1180
<< nsubdiffcont >>
rect -100 640 -80 765
rect 1000 640 1020 765
rect -100 95 -80 365
rect 1000 95 1020 365
rect -100 -795 -80 -225
rect 1000 -795 1020 -225
<< poly >>
rect -15 775 35 790
rect 85 775 135 790
rect 185 775 235 790
rect 285 775 335 790
rect 385 775 435 790
rect 485 775 535 790
rect 585 775 635 790
rect 685 775 735 790
rect 785 775 835 790
rect 885 775 935 790
rect -15 610 35 625
rect 85 615 135 625
rect 185 615 235 625
rect 285 615 335 625
rect 385 615 435 625
rect 485 615 535 625
rect 585 615 635 625
rect 685 615 735 625
rect 785 615 835 625
rect -60 600 35 610
rect -60 580 -50 600
rect -30 595 35 600
rect 60 600 835 615
rect 885 610 935 625
rect 885 600 980 610
rect -30 580 -20 595
rect -60 570 -20 580
rect 60 545 75 600
rect 885 595 950 600
rect 940 580 950 595
rect 970 580 980 600
rect 940 570 980 580
rect -60 535 75 545
rect -60 515 -50 535
rect -30 530 75 535
rect -30 515 -20 530
rect -60 505 -20 515
rect 0 475 40 485
rect 0 455 10 475
rect 30 460 40 475
rect 95 460 135 465
rect 30 455 135 460
rect 0 445 135 455
rect 85 435 135 445
rect -60 425 -20 435
rect -60 405 -50 425
rect -30 410 -20 425
rect 85 420 835 435
rect -30 405 35 410
rect -60 395 35 405
rect -15 380 35 395
rect 85 380 135 420
rect 185 380 235 395
rect 285 380 335 395
rect 385 380 435 420
rect 485 380 535 420
rect 585 380 635 395
rect 685 380 735 395
rect 785 380 835 420
rect 940 425 980 435
rect 940 410 950 425
rect 885 405 950 410
rect 970 405 980 425
rect 885 395 980 405
rect 885 380 935 395
rect -15 65 35 80
rect 85 65 135 80
rect 185 40 235 80
rect 285 40 335 80
rect 385 65 435 80
rect 485 65 535 80
rect 585 40 635 80
rect 685 40 735 80
rect 785 65 835 80
rect 885 65 935 80
rect -5 30 735 40
rect -5 10 5 30
rect 25 25 735 30
rect 25 10 35 25
rect -5 0 35 10
rect 240 -10 280 0
rect 240 -30 250 -10
rect 270 -25 280 -10
rect 640 -10 680 0
rect 640 -25 650 -10
rect 270 -30 650 -25
rect 670 -30 680 -10
rect 240 -40 680 -30
rect -5 -110 35 -100
rect -5 -130 5 -110
rect 25 -125 35 -110
rect 25 -130 835 -125
rect -5 -140 835 -130
rect -60 -165 -20 -155
rect -60 -185 -50 -165
rect -30 -180 -20 -165
rect -30 -185 35 -180
rect -60 -195 35 -185
rect -15 -210 35 -195
rect 85 -210 135 -140
rect 185 -210 235 -195
rect 285 -210 335 -195
rect 385 -210 435 -140
rect 485 -210 535 -140
rect 585 -210 635 -195
rect 685 -210 735 -195
rect 785 -210 835 -140
rect 940 -165 980 -155
rect 940 -180 950 -165
rect 885 -185 950 -180
rect 970 -185 980 -165
rect 885 -195 980 -185
rect 885 -210 935 -195
rect -15 -825 35 -810
rect 85 -825 135 -810
rect 185 -850 235 -810
rect 285 -850 335 -810
rect 385 -825 435 -810
rect 485 -825 535 -810
rect 585 -850 635 -810
rect 685 -850 735 -810
rect 785 -825 835 -810
rect 885 -825 935 -810
rect 185 -860 735 -850
rect 185 -865 450 -860
rect 440 -880 450 -865
rect 470 -865 735 -860
rect 470 -880 480 -865
rect 440 -890 480 -880
rect 450 -950 470 -890
rect 380 -960 540 -950
rect 380 -980 390 -960
rect 410 -965 510 -960
rect 410 -980 420 -965
rect 380 -990 420 -980
rect 500 -980 510 -965
rect 530 -980 540 -960
rect 500 -990 540 -980
rect -60 -1060 -20 -1050
rect -60 -1080 -50 -1060
rect -30 -1075 -20 -1060
rect -30 -1080 100 -1075
rect -60 -1090 100 -1080
rect 85 -1110 100 -1090
rect -60 -1125 -20 -1115
rect -60 -1145 -50 -1125
rect -30 -1140 -20 -1125
rect 85 -1125 835 -1110
rect -30 -1145 35 -1140
rect -60 -1155 35 -1145
rect -15 -1165 35 -1155
rect 85 -1165 135 -1125
rect 185 -1165 235 -1150
rect 285 -1165 335 -1150
rect 385 -1165 435 -1125
rect 485 -1165 535 -1125
rect 585 -1165 635 -1150
rect 685 -1165 735 -1150
rect 785 -1165 835 -1125
rect 940 -1125 980 -1115
rect 940 -1140 950 -1125
rect 885 -1145 950 -1140
rect 970 -1145 980 -1125
rect 885 -1155 980 -1145
rect 885 -1165 935 -1155
rect -15 -1780 35 -1765
rect 85 -1780 135 -1765
rect 185 -1800 235 -1765
rect 285 -1800 335 -1765
rect 385 -1780 435 -1765
rect 485 -1780 535 -1765
rect -65 -1805 -25 -1800
rect 185 -1805 335 -1800
rect 585 -1805 635 -1765
rect 685 -1805 735 -1765
rect 785 -1780 835 -1765
rect 885 -1780 935 -1765
rect -65 -1810 735 -1805
rect -65 -1830 -55 -1810
rect -35 -1820 735 -1810
rect -35 -1830 -25 -1820
rect -65 -1840 -25 -1830
<< polycont >>
rect -50 580 -30 600
rect 950 580 970 600
rect -50 515 -30 535
rect 10 455 30 475
rect -50 405 -30 425
rect 950 405 970 425
rect 5 10 25 30
rect 250 -30 270 -10
rect 650 -30 670 -10
rect 5 -130 25 -110
rect -50 -185 -30 -165
rect 950 -185 970 -165
rect 450 -880 470 -860
rect 390 -980 410 -960
rect 510 -980 530 -960
rect -50 -1080 -30 -1060
rect -50 -1145 -30 -1125
rect 950 -1145 970 -1125
rect -55 -1830 -35 -1810
<< locali >>
rect -110 765 -20 770
rect -110 640 -100 765
rect -80 640 -50 765
rect -30 640 -20 765
rect -110 630 -20 640
rect 40 765 80 770
rect 40 640 50 765
rect 70 640 80 765
rect 40 630 80 640
rect 140 765 180 770
rect 140 640 150 765
rect 170 640 180 765
rect -60 600 -20 630
rect -60 580 -50 600
rect -30 580 -20 600
rect -60 570 -20 580
rect 140 610 180 640
rect 240 765 280 770
rect 240 640 250 765
rect 270 640 280 765
rect 240 630 280 640
rect 340 765 380 770
rect 340 640 350 765
rect 370 640 380 765
rect 340 610 380 640
rect 440 765 480 770
rect 440 640 450 765
rect 470 640 480 765
rect 440 630 480 640
rect 540 765 580 770
rect 540 640 550 765
rect 570 640 580 765
rect 540 610 580 640
rect 640 765 680 770
rect 640 640 650 765
rect 670 640 680 765
rect 640 630 680 640
rect 740 765 780 770
rect 740 640 750 765
rect 770 640 780 765
rect 740 610 780 640
rect 840 765 880 770
rect 840 640 850 765
rect 870 640 880 765
rect 840 630 880 640
rect 940 765 1030 770
rect 940 640 950 765
rect 970 640 1000 765
rect 1020 640 1030 765
rect 940 630 1030 640
rect 140 590 780 610
rect -115 535 -20 545
rect -115 525 -50 535
rect -60 515 -50 525
rect -30 515 -20 535
rect -60 505 -20 515
rect -115 475 40 485
rect -115 465 10 475
rect 0 455 10 465
rect 30 455 40 475
rect 0 445 40 455
rect -60 425 -20 435
rect -60 405 -50 425
rect -30 405 -20 425
rect -60 375 -20 405
rect -110 365 -20 375
rect -110 95 -100 365
rect -80 95 -50 365
rect -30 95 -20 365
rect -110 85 -20 95
rect 40 365 80 375
rect 40 95 50 365
rect 70 95 80 365
rect 40 85 80 95
rect 140 365 180 590
rect 140 95 150 365
rect 170 95 180 365
rect 140 85 180 95
rect 240 365 280 375
rect 240 95 250 365
rect 270 95 280 365
rect -120 30 35 40
rect -120 20 5 30
rect -5 10 5 20
rect 25 10 35 30
rect -5 0 35 10
rect 60 -40 80 85
rect 240 -10 280 95
rect 340 365 380 590
rect 340 95 350 365
rect 370 95 380 365
rect 340 85 380 95
rect 440 365 480 375
rect 440 95 450 365
rect 470 95 480 365
rect 440 85 480 95
rect 540 365 580 590
rect 540 95 550 365
rect 570 95 580 365
rect 540 85 580 95
rect 640 365 680 375
rect 640 95 650 365
rect 670 95 680 365
rect 240 -30 250 -10
rect 270 -30 280 -10
rect 240 -40 280 -30
rect 60 -50 100 -40
rect 60 -70 70 -50
rect 90 -60 100 -50
rect 450 -60 470 85
rect 640 -10 680 95
rect 740 365 780 590
rect 940 600 980 630
rect 940 580 950 600
rect 970 580 980 600
rect 940 570 980 580
rect 940 425 980 435
rect 940 405 950 425
rect 970 405 980 425
rect 940 375 980 405
rect 740 95 750 365
rect 770 95 780 365
rect 740 85 780 95
rect 840 365 880 375
rect 840 95 850 365
rect 870 95 880 365
rect 840 85 880 95
rect 940 365 1030 375
rect 940 95 950 365
rect 970 95 1000 365
rect 1020 95 1030 365
rect 940 85 1030 95
rect 640 -30 650 -10
rect 670 -30 680 -10
rect 640 -40 680 -30
rect 840 -60 860 85
rect 90 -70 860 -60
rect 60 -80 860 -70
rect -120 -110 35 -100
rect -120 -120 5 -110
rect -5 -130 5 -120
rect 25 -130 35 -110
rect -5 -140 35 -130
rect 140 -155 780 -135
rect -60 -165 -20 -155
rect -60 -185 -50 -165
rect -30 -185 -20 -165
rect -60 -215 -20 -185
rect -110 -225 -20 -215
rect -110 -795 -100 -225
rect -80 -795 -50 -225
rect -30 -795 -20 -225
rect -110 -805 -20 -795
rect 40 -225 80 -215
rect 40 -795 50 -225
rect 70 -795 80 -225
rect 40 -910 80 -795
rect 140 -225 180 -155
rect 340 -195 580 -175
rect 140 -795 150 -225
rect 170 -795 180 -225
rect 140 -805 180 -795
rect 240 -225 280 -215
rect 240 -795 250 -225
rect 270 -795 280 -225
rect 240 -805 280 -795
rect 340 -225 380 -195
rect 340 -795 350 -225
rect 370 -795 380 -225
rect 340 -805 380 -795
rect 440 -225 480 -215
rect 440 -795 450 -225
rect 470 -795 480 -225
rect 440 -860 480 -795
rect 540 -225 580 -195
rect 540 -795 550 -225
rect 570 -795 580 -225
rect 540 -805 580 -795
rect 640 -225 680 -215
rect 640 -795 650 -225
rect 670 -795 680 -225
rect 640 -805 680 -795
rect 740 -225 780 -155
rect 940 -165 980 -155
rect 940 -185 950 -165
rect 970 -185 980 -165
rect 940 -215 980 -185
rect 740 -795 750 -225
rect 770 -795 780 -225
rect 740 -805 780 -795
rect 840 -225 880 -215
rect 840 -795 850 -225
rect 870 -795 880 -225
rect 440 -880 450 -860
rect 470 -880 480 -860
rect 440 -890 480 -880
rect 840 -910 880 -795
rect 940 -225 1030 -215
rect 940 -795 950 -225
rect 970 -795 1000 -225
rect 1020 -795 1030 -225
rect 940 -805 1030 -795
rect 40 -930 1035 -910
rect 40 -960 420 -950
rect 40 -970 390 -960
rect -60 -1060 -20 -1050
rect -60 -1070 -50 -1060
rect -115 -1080 -50 -1070
rect -30 -1080 -20 -1060
rect -115 -1090 -20 -1080
rect -60 -1125 -20 -1115
rect -60 -1145 -50 -1125
rect -30 -1145 -20 -1125
rect -60 -1170 -20 -1145
rect -110 -1180 -20 -1170
rect -110 -1750 -100 -1180
rect -80 -1750 -50 -1180
rect -30 -1750 -20 -1180
rect -110 -1760 -20 -1750
rect 40 -1180 80 -970
rect 380 -980 390 -970
rect 410 -980 420 -960
rect 380 -990 420 -980
rect 40 -1750 50 -1180
rect 70 -1750 80 -1180
rect 40 -1760 80 -1750
rect 140 -1000 180 -990
rect 140 -1020 150 -1000
rect 170 -1020 180 -1000
rect 140 -1180 180 -1020
rect 140 -1750 150 -1180
rect 170 -1750 180 -1180
rect -115 -1810 -25 -1800
rect -115 -1820 -55 -1810
rect -65 -1830 -55 -1820
rect -35 -1830 -25 -1810
rect -65 -1840 -25 -1830
rect 140 -1820 180 -1750
rect 240 -1180 280 -1170
rect 240 -1750 250 -1180
rect 270 -1750 280 -1180
rect 240 -1760 280 -1750
rect 340 -1180 380 -1170
rect 340 -1750 350 -1180
rect 370 -1750 380 -1180
rect 340 -1780 380 -1750
rect 440 -1180 480 -930
rect 500 -960 880 -950
rect 500 -980 510 -960
rect 530 -970 880 -960
rect 530 -980 540 -970
rect 500 -990 540 -980
rect 440 -1750 450 -1180
rect 470 -1750 480 -1180
rect 440 -1760 480 -1750
rect 540 -1045 580 -1035
rect 540 -1065 550 -1045
rect 570 -1065 580 -1045
rect 540 -1180 580 -1065
rect 540 -1750 550 -1180
rect 570 -1750 580 -1180
rect 540 -1780 580 -1750
rect 640 -1180 680 -1170
rect 640 -1750 650 -1180
rect 670 -1750 680 -1180
rect 640 -1760 680 -1750
rect 740 -1180 780 -1170
rect 740 -1750 750 -1180
rect 770 -1750 780 -1180
rect 340 -1800 580 -1780
rect 740 -1820 780 -1750
rect 840 -1180 880 -970
rect 840 -1750 850 -1180
rect 870 -1750 880 -1180
rect 840 -1760 880 -1750
rect 940 -1125 980 -1115
rect 940 -1145 950 -1125
rect 970 -1145 980 -1125
rect 940 -1170 980 -1145
rect 940 -1180 1030 -1170
rect 940 -1750 950 -1180
rect 970 -1750 1000 -1180
rect 1020 -1750 1030 -1180
rect 940 -1760 1030 -1750
rect 140 -1840 780 -1820
<< viali >>
rect -100 640 -80 765
rect -50 640 -30 765
rect 50 640 70 765
rect 250 640 270 765
rect 450 640 470 765
rect 650 640 670 765
rect 850 640 870 765
rect 950 640 970 765
rect 1000 640 1020 765
rect -100 95 -80 365
rect -50 95 -30 365
rect 70 -70 90 -50
rect 950 95 970 365
rect 1000 95 1020 365
rect 650 -30 670 -10
rect -100 -795 -80 -225
rect -50 -795 -30 -225
rect 250 -795 270 -225
rect 650 -795 670 -225
rect 950 -795 970 -225
rect 1000 -795 1020 -225
rect -100 -1750 -80 -1180
rect -50 -1750 -30 -1180
rect 150 -1020 170 -1000
rect 250 -1750 270 -1180
rect 550 -1065 570 -1045
rect 650 -1750 670 -1180
rect 950 -1750 970 -1180
rect 1000 -1750 1020 -1180
<< metal1 >>
rect -115 765 1035 770
rect -115 640 -100 765
rect -80 640 -50 765
rect -30 640 50 765
rect 70 640 250 765
rect 270 640 450 765
rect 470 640 650 765
rect 670 640 850 765
rect 870 640 950 765
rect 970 640 1000 765
rect 1020 640 1035 765
rect -115 365 1035 640
rect -115 95 -100 365
rect -80 95 -50 365
rect -30 95 950 365
rect 970 95 1000 365
rect 1020 95 1035 365
rect -115 85 1035 95
rect -115 -215 -15 85
rect 540 -10 680 0
rect 540 -30 650 -10
rect 670 -30 680 -10
rect 540 -40 680 -30
rect 60 -50 380 -40
rect 60 -70 70 -50
rect 90 -70 380 -50
rect 60 -80 380 -70
rect -115 -225 280 -215
rect -115 -795 -100 -225
rect -80 -795 -50 -225
rect -30 -795 250 -225
rect 270 -795 280 -225
rect -115 -805 280 -795
rect 340 -990 380 -80
rect 140 -1000 380 -990
rect 140 -1020 150 -1000
rect 170 -1020 380 -1000
rect 140 -1030 380 -1020
rect 540 -1045 580 -40
rect 935 -215 1035 85
rect 640 -225 1035 -215
rect 640 -795 650 -225
rect 670 -795 950 -225
rect 970 -795 1000 -225
rect 1020 -795 1035 -225
rect 640 -805 1035 -795
rect 540 -1065 550 -1045
rect 570 -1065 580 -1045
rect 540 -1075 580 -1065
rect -115 -1180 1035 -1170
rect -115 -1750 -100 -1180
rect -80 -1750 -50 -1180
rect -30 -1750 250 -1180
rect 270 -1750 650 -1180
rect 670 -1750 950 -1180
rect 970 -1750 1000 -1180
rect 1020 -1750 1035 -1180
rect -115 -1760 1035 -1750
<< labels >>
rlabel locali 1035 -920 1035 -920 3 Vout
rlabel metal1 -115 700 -115 700 7 Vp
rlabel locali -115 535 -115 535 7 Vbp
rlabel locali -115 475 -115 475 7 V1
rlabel locali -120 30 -120 30 7 V2
rlabel locali -120 -110 -120 -110 7 Vcp
rlabel locali -115 -1080 -115 -1080 7 Vcn
rlabel locali -115 -1810 -115 -1810 7 Vbn
rlabel metal1 -115 -1470 -115 -1470 7 Vn
<< end >>
