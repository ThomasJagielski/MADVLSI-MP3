magic
tech sky130A
timestamp 1615701304
<< locali >>
rect 1330 3270 1360 3290
rect 2490 2975 2510 2995
rect 20 2525 40 2565
rect 2490 2535 2510 2555
rect 1330 1640 1360 1660
rect 1330 1560 1360 1580
rect 2490 1565 2510 1585
rect 1325 0 1365 20
<< metal1 >>
rect 20 2645 45 3240
rect 1325 1720 1360 3240
rect 20 60 45 650
rect 1325 60 1365 650
use differential_pair  differential_pair_0
timestamp 1615700760
transform 1 0 1475 0 1 2520
box -135 -2540 1055 780
use cascode_bias  cascode_bias_0
timestamp 1615699134
transform 1 0 120 0 1 2630
box -120 -2630 1230 670
<< labels >>
rlabel metal1 20 2945 20 2945 7 VP
rlabel locali 20 2545 20 2545 7 Vbp
rlabel metal1 20 355 20 355 7 VN
rlabel locali 2510 1575 2510 1575 3 Vout
rlabel locali 2510 2985 2510 2985 3 V1
rlabel locali 2490 2535 2510 2555 3 V2
<< end >>
