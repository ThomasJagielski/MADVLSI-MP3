magic
tech sky130A
timestamp 1615644373
<< nmos >>
rect 0 0 50 600
rect 100 0 150 600
rect 200 0 250 600
rect 380 0 430 600
rect 480 0 530 600
rect 580 0 630 600
rect 680 0 730 600
rect 860 0 910 600
rect 960 0 1010 600
rect 1060 0 1110 600
rect 0 -1000 50 -400
rect 100 -1000 150 -400
rect 200 -1000 250 -400
rect 300 -1000 350 -400
rect 480 -1000 530 -400
rect 580 -1000 630 -400
rect 760 -1000 810 -400
rect 860 -1000 910 -400
rect 960 -1000 1010 -400
rect 1060 -1000 1110 -400
rect 0 -2000 50 -1400
rect 100 -2000 150 -1400
rect 200 -2000 250 -1400
rect 300 -2000 350 -1400
rect 480 -2000 530 -1400
rect 580 -2000 630 -1400
rect 760 -2000 810 -1400
rect 860 -2000 910 -1400
rect 960 -2000 1010 -1400
rect 1060 -2000 1110 -1400
rect 0 -3000 50 -2400
rect 100 -3000 150 -2400
rect 200 -3000 250 -2400
rect 300 -3000 350 -2400
rect 480 -3000 530 -2400
rect 580 -3000 630 -2400
rect 760 -3000 810 -2400
rect 860 -3000 910 -2400
rect 960 -3000 1010 -2400
rect 1060 -3000 1110 -2400
<< ndiff >>
rect -50 585 0 600
rect -50 15 -35 585
rect -15 15 0 585
rect -50 0 0 15
rect 50 585 100 600
rect 50 15 65 585
rect 85 15 100 585
rect 50 0 100 15
rect 150 585 200 600
rect 150 15 165 585
rect 185 15 200 585
rect 150 0 200 15
rect 250 585 300 600
rect 250 15 265 585
rect 285 15 300 585
rect 250 0 300 15
rect 330 585 380 600
rect 330 15 345 585
rect 365 15 380 585
rect 330 0 380 15
rect 430 585 480 600
rect 430 15 445 585
rect 465 15 480 585
rect 430 0 480 15
rect 530 585 580 600
rect 530 15 545 585
rect 565 15 580 585
rect 530 0 580 15
rect 630 585 680 600
rect 630 15 645 585
rect 665 15 680 585
rect 630 0 680 15
rect 730 585 780 600
rect 730 15 745 585
rect 765 15 780 585
rect 730 0 780 15
rect 810 585 860 600
rect 810 15 825 585
rect 845 15 860 585
rect 810 0 860 15
rect 910 585 960 600
rect 910 15 925 585
rect 945 15 960 585
rect 910 0 960 15
rect 1010 585 1060 600
rect 1010 15 1025 585
rect 1045 15 1060 585
rect 1010 0 1060 15
rect 1110 585 1160 600
rect 1110 15 1125 585
rect 1145 15 1160 585
rect 1110 0 1160 15
rect -50 -415 0 -400
rect -50 -985 -35 -415
rect -15 -985 0 -415
rect -50 -1000 0 -985
rect 50 -415 100 -400
rect 50 -985 65 -415
rect 85 -985 100 -415
rect 50 -1000 100 -985
rect 150 -415 200 -400
rect 150 -985 165 -415
rect 185 -985 200 -415
rect 150 -1000 200 -985
rect 250 -415 300 -400
rect 250 -985 265 -415
rect 285 -985 300 -415
rect 250 -1000 300 -985
rect 350 -415 400 -400
rect 350 -985 365 -415
rect 385 -985 400 -415
rect 350 -1000 400 -985
rect 430 -415 480 -400
rect 430 -985 445 -415
rect 465 -985 480 -415
rect 430 -1000 480 -985
rect 530 -415 580 -400
rect 530 -985 545 -415
rect 565 -985 580 -415
rect 530 -1000 580 -985
rect 630 -415 680 -400
rect 630 -985 645 -415
rect 665 -985 680 -415
rect 630 -1000 680 -985
rect 710 -415 760 -400
rect 710 -985 725 -415
rect 745 -985 760 -415
rect 710 -1000 760 -985
rect 810 -415 860 -400
rect 810 -985 825 -415
rect 845 -985 860 -415
rect 810 -1000 860 -985
rect 910 -415 960 -400
rect 910 -985 925 -415
rect 945 -985 960 -415
rect 910 -1000 960 -985
rect 1010 -415 1060 -400
rect 1010 -985 1025 -415
rect 1045 -985 1060 -415
rect 1010 -1000 1060 -985
rect 1110 -415 1160 -400
rect 1110 -985 1125 -415
rect 1145 -985 1160 -415
rect 1110 -1000 1160 -985
rect -50 -1415 0 -1400
rect -50 -1985 -35 -1415
rect -15 -1985 0 -1415
rect -50 -2000 0 -1985
rect 50 -1415 100 -1400
rect 50 -1985 65 -1415
rect 85 -1985 100 -1415
rect 50 -2000 100 -1985
rect 150 -1415 200 -1400
rect 150 -1985 165 -1415
rect 185 -1985 200 -1415
rect 150 -2000 200 -1985
rect 250 -1415 300 -1400
rect 250 -1985 265 -1415
rect 285 -1985 300 -1415
rect 250 -2000 300 -1985
rect 350 -1415 400 -1400
rect 350 -1985 365 -1415
rect 385 -1985 400 -1415
rect 350 -2000 400 -1985
rect 430 -1415 480 -1400
rect 430 -1985 445 -1415
rect 465 -1985 480 -1415
rect 430 -2000 480 -1985
rect 530 -1415 580 -1400
rect 530 -1985 545 -1415
rect 565 -1985 580 -1415
rect 530 -2000 580 -1985
rect 630 -1415 680 -1400
rect 630 -1985 645 -1415
rect 665 -1985 680 -1415
rect 630 -2000 680 -1985
rect 710 -1415 760 -1400
rect 710 -1985 725 -1415
rect 745 -1985 760 -1415
rect 710 -2000 760 -1985
rect 810 -1415 860 -1400
rect 810 -1985 825 -1415
rect 845 -1985 860 -1415
rect 810 -2000 860 -1985
rect 910 -1415 960 -1400
rect 910 -1985 925 -1415
rect 945 -1985 960 -1415
rect 910 -2000 960 -1985
rect 1010 -1415 1060 -1400
rect 1010 -1985 1025 -1415
rect 1045 -1985 1060 -1415
rect 1010 -2000 1060 -1985
rect 1110 -1415 1160 -1400
rect 1110 -1985 1125 -1415
rect 1145 -1985 1160 -1415
rect 1110 -2000 1160 -1985
rect -50 -2415 0 -2400
rect -50 -2985 -35 -2415
rect -15 -2985 0 -2415
rect -50 -3000 0 -2985
rect 50 -2415 100 -2400
rect 50 -2985 65 -2415
rect 85 -2985 100 -2415
rect 50 -3000 100 -2985
rect 150 -2415 200 -2400
rect 150 -2985 165 -2415
rect 185 -2985 200 -2415
rect 150 -3000 200 -2985
rect 250 -2415 300 -2400
rect 250 -2985 265 -2415
rect 285 -2985 300 -2415
rect 250 -3000 300 -2985
rect 350 -2415 400 -2400
rect 350 -2985 365 -2415
rect 385 -2985 400 -2415
rect 350 -3000 400 -2985
rect 430 -2415 480 -2400
rect 430 -2985 445 -2415
rect 465 -2985 480 -2415
rect 430 -3000 480 -2985
rect 530 -2415 580 -2400
rect 530 -2985 545 -2415
rect 565 -2985 580 -2415
rect 530 -3000 580 -2985
rect 630 -2415 680 -2400
rect 630 -2985 645 -2415
rect 665 -2985 680 -2415
rect 630 -3000 680 -2985
rect 710 -2415 760 -2400
rect 710 -2985 725 -2415
rect 745 -2985 760 -2415
rect 710 -3000 760 -2985
rect 810 -2415 860 -2400
rect 810 -2985 825 -2415
rect 845 -2985 860 -2415
rect 810 -3000 860 -2985
rect 910 -2415 960 -2400
rect 910 -2985 925 -2415
rect 945 -2985 960 -2415
rect 910 -3000 960 -2985
rect 1010 -2415 1060 -2400
rect 1010 -2985 1025 -2415
rect 1045 -2985 1060 -2415
rect 1010 -3000 1060 -2985
rect 1110 -2415 1160 -2400
rect 1110 -2985 1125 -2415
rect 1145 -2985 1160 -2415
rect 1110 -3000 1160 -2985
<< ndiffc >>
rect -35 15 -15 585
rect 65 15 85 585
rect 165 15 185 585
rect 265 15 285 585
rect 345 15 365 585
rect 445 15 465 585
rect 545 15 565 585
rect 645 15 665 585
rect 745 15 765 585
rect 825 15 845 585
rect 925 15 945 585
rect 1025 15 1045 585
rect 1125 15 1145 585
rect -35 -985 -15 -415
rect 65 -985 85 -415
rect 165 -985 185 -415
rect 265 -985 285 -415
rect 365 -985 385 -415
rect 445 -985 465 -415
rect 545 -985 565 -415
rect 645 -985 665 -415
rect 725 -985 745 -415
rect 825 -985 845 -415
rect 925 -985 945 -415
rect 1025 -985 1045 -415
rect 1125 -985 1145 -415
rect -35 -1985 -15 -1415
rect 65 -1985 85 -1415
rect 165 -1985 185 -1415
rect 265 -1985 285 -1415
rect 365 -1985 385 -1415
rect 445 -1985 465 -1415
rect 545 -1985 565 -1415
rect 645 -1985 665 -1415
rect 725 -1985 745 -1415
rect 825 -1985 845 -1415
rect 925 -1985 945 -1415
rect 1025 -1985 1045 -1415
rect 1125 -1985 1145 -1415
rect -35 -2985 -15 -2415
rect 65 -2985 85 -2415
rect 165 -2985 185 -2415
rect 265 -2985 285 -2415
rect 365 -2985 385 -2415
rect 445 -2985 465 -2415
rect 545 -2985 565 -2415
rect 645 -2985 665 -2415
rect 725 -2985 745 -2415
rect 825 -2985 845 -2415
rect 925 -2985 945 -2415
rect 1025 -2985 1045 -2415
rect 1125 -2985 1145 -2415
<< psubdiff >>
rect -100 585 -50 600
rect -100 15 -85 585
rect -65 15 -50 585
rect -100 0 -50 15
rect 1160 585 1210 600
rect 1160 15 1175 585
rect 1195 15 1210 585
rect 1160 0 1210 15
rect -100 -415 -50 -400
rect -100 -985 -85 -415
rect -65 -985 -50 -415
rect -100 -1000 -50 -985
rect 1160 -415 1210 -400
rect 1160 -985 1175 -415
rect 1195 -985 1210 -415
rect 1160 -1000 1210 -985
rect -100 -1415 -50 -1400
rect -100 -1985 -85 -1415
rect -65 -1985 -50 -1415
rect -100 -2000 -50 -1985
rect 1160 -1415 1210 -1400
rect 1160 -1985 1175 -1415
rect 1195 -1985 1210 -1415
rect 1160 -2000 1210 -1985
rect -100 -2415 -50 -2400
rect -100 -2985 -85 -2415
rect -65 -2985 -50 -2415
rect -100 -3000 -50 -2985
rect 1160 -2415 1210 -2400
rect 1160 -2985 1175 -2415
rect 1195 -2985 1210 -2415
rect 1160 -3000 1210 -2985
<< psubdiffcont >>
rect -85 15 -65 585
rect 1175 15 1195 585
rect -85 -985 -65 -415
rect 1175 -985 1195 -415
rect -85 -1985 -65 -1415
rect 1175 -1985 1195 -1415
rect -85 -2985 -65 -2415
rect 1175 -2985 1195 -2415
<< poly >>
rect 0 600 50 615
rect 100 600 150 615
rect 200 600 250 615
rect 380 600 430 615
rect 480 600 530 615
rect 580 600 630 615
rect 680 600 730 615
rect 860 600 910 615
rect 960 600 1010 615
rect 1060 600 1110 615
rect 0 -15 50 0
rect 100 -15 150 0
rect 200 -15 250 0
rect 380 -15 430 0
rect 480 -15 530 0
rect 580 -15 630 0
rect 680 -15 730 0
rect 860 -15 910 0
rect 960 -15 1010 0
rect 1060 -15 1110 0
rect 0 -400 50 -385
rect 100 -400 150 -385
rect 200 -400 250 -385
rect 300 -400 350 -385
rect 480 -400 530 -385
rect 580 -400 630 -385
rect 760 -400 810 -385
rect 860 -400 910 -385
rect 960 -400 1010 -385
rect 1060 -400 1110 -385
rect 0 -1015 50 -1000
rect 100 -1015 150 -1000
rect 200 -1015 250 -1000
rect 300 -1015 350 -1000
rect 480 -1015 530 -1000
rect 580 -1015 630 -1000
rect 760 -1015 810 -1000
rect 860 -1015 910 -1000
rect 960 -1015 1010 -1000
rect 1060 -1015 1110 -1000
rect 0 -1400 50 -1385
rect 100 -1400 150 -1385
rect 200 -1400 250 -1385
rect 300 -1400 350 -1385
rect 480 -1400 530 -1385
rect 580 -1400 630 -1385
rect 760 -1400 810 -1385
rect 860 -1400 910 -1385
rect 960 -1400 1010 -1385
rect 1060 -1400 1110 -1385
rect 0 -2015 50 -2000
rect 100 -2015 150 -2000
rect 200 -2015 250 -2000
rect 300 -2015 350 -2000
rect 480 -2015 530 -2000
rect 580 -2015 630 -2000
rect 760 -2015 810 -2000
rect 860 -2015 910 -2000
rect 960 -2015 1010 -2000
rect 1060 -2015 1110 -2000
rect 0 -2400 50 -2385
rect 100 -2400 150 -2385
rect 200 -2400 250 -2385
rect 300 -2400 350 -2385
rect 480 -2400 530 -2385
rect 580 -2400 630 -2385
rect 760 -2400 810 -2385
rect 860 -2400 910 -2385
rect 960 -2400 1010 -2385
rect 1060 -2400 1110 -2385
rect 0 -3015 50 -3000
rect 100 -3015 150 -3000
rect 200 -3015 250 -3000
rect 300 -3015 350 -3000
rect 480 -3015 530 -3000
rect 580 -3015 630 -3000
rect 760 -3015 810 -3000
rect 860 -3015 910 -3000
rect 960 -3015 1010 -3000
rect 1060 -3015 1110 -3000
<< locali >>
rect -95 585 -5 595
rect -95 15 -85 585
rect -65 15 -35 585
rect -15 15 -5 585
rect -95 5 -5 15
rect 55 585 95 595
rect 55 15 65 585
rect 85 15 95 585
rect 55 5 95 15
rect 155 585 195 595
rect 155 15 165 585
rect 185 15 195 585
rect 155 5 195 15
rect 255 585 295 595
rect 255 15 265 585
rect 285 15 295 585
rect 255 5 295 15
rect 335 585 375 595
rect 335 15 345 585
rect 365 15 375 585
rect 335 5 375 15
rect 435 585 475 595
rect 435 15 445 585
rect 465 15 475 585
rect 435 5 475 15
rect 535 585 575 595
rect 535 15 545 585
rect 565 15 575 585
rect 535 5 575 15
rect 635 585 675 595
rect 635 15 645 585
rect 665 15 675 585
rect 635 5 675 15
rect 735 585 775 595
rect 735 15 745 585
rect 765 15 775 585
rect 735 5 775 15
rect 815 585 855 595
rect 815 15 825 585
rect 845 15 855 585
rect 815 5 855 15
rect 915 585 955 595
rect 915 15 925 585
rect 945 15 955 585
rect 915 5 955 15
rect 1015 585 1055 595
rect 1015 15 1025 585
rect 1045 15 1055 585
rect 1015 5 1055 15
rect 1115 585 1205 595
rect 1115 15 1125 585
rect 1145 15 1175 585
rect 1195 15 1205 585
rect 1115 5 1205 15
rect -95 -415 -5 -405
rect -95 -985 -85 -415
rect -65 -985 -35 -415
rect -15 -985 -5 -415
rect -95 -995 -5 -985
rect 55 -415 95 -405
rect 55 -985 65 -415
rect 85 -985 95 -415
rect 55 -995 95 -985
rect 155 -415 195 -405
rect 155 -985 165 -415
rect 185 -985 195 -415
rect 155 -995 195 -985
rect 255 -415 295 -405
rect 255 -985 265 -415
rect 285 -985 295 -415
rect 255 -995 295 -985
rect 355 -415 395 -405
rect 355 -985 365 -415
rect 385 -985 395 -415
rect 355 -995 395 -985
rect 435 -415 475 -405
rect 435 -985 445 -415
rect 465 -985 475 -415
rect 435 -995 475 -985
rect 535 -415 575 -405
rect 535 -985 545 -415
rect 565 -985 575 -415
rect 535 -995 575 -985
rect 635 -415 675 -405
rect 635 -985 645 -415
rect 665 -985 675 -415
rect 635 -995 675 -985
rect 715 -415 755 -405
rect 715 -985 725 -415
rect 745 -985 755 -415
rect 715 -995 755 -985
rect 815 -415 855 -405
rect 815 -985 825 -415
rect 845 -985 855 -415
rect 815 -995 855 -985
rect 915 -415 955 -405
rect 915 -985 925 -415
rect 945 -985 955 -415
rect 915 -995 955 -985
rect 1015 -415 1055 -405
rect 1015 -985 1025 -415
rect 1045 -985 1055 -415
rect 1015 -995 1055 -985
rect 1115 -415 1205 -405
rect 1115 -985 1125 -415
rect 1145 -985 1175 -415
rect 1195 -985 1205 -415
rect 1115 -995 1205 -985
rect -95 -1415 -5 -1405
rect -95 -1985 -85 -1415
rect -65 -1985 -35 -1415
rect -15 -1985 -5 -1415
rect -95 -1995 -5 -1985
rect 55 -1415 95 -1405
rect 55 -1985 65 -1415
rect 85 -1985 95 -1415
rect 55 -1995 95 -1985
rect 155 -1415 195 -1405
rect 155 -1985 165 -1415
rect 185 -1985 195 -1415
rect 155 -1995 195 -1985
rect 255 -1415 295 -1405
rect 255 -1985 265 -1415
rect 285 -1985 295 -1415
rect 255 -1995 295 -1985
rect 355 -1415 395 -1405
rect 355 -1985 365 -1415
rect 385 -1985 395 -1415
rect 355 -1995 395 -1985
rect 435 -1415 475 -1405
rect 435 -1985 445 -1415
rect 465 -1985 475 -1415
rect 435 -1995 475 -1985
rect 535 -1415 575 -1405
rect 535 -1985 545 -1415
rect 565 -1985 575 -1415
rect 535 -1995 575 -1985
rect 635 -1415 675 -1405
rect 635 -1985 645 -1415
rect 665 -1985 675 -1415
rect 635 -1995 675 -1985
rect 715 -1415 755 -1405
rect 715 -1985 725 -1415
rect 745 -1985 755 -1415
rect 715 -1995 755 -1985
rect 815 -1415 855 -1405
rect 815 -1985 825 -1415
rect 845 -1985 855 -1415
rect 815 -1995 855 -1985
rect 915 -1415 955 -1405
rect 915 -1985 925 -1415
rect 945 -1985 955 -1415
rect 915 -1995 955 -1985
rect 1015 -1415 1055 -1405
rect 1015 -1985 1025 -1415
rect 1045 -1985 1055 -1415
rect 1015 -1995 1055 -1985
rect 1115 -1415 1205 -1405
rect 1115 -1985 1125 -1415
rect 1145 -1985 1175 -1415
rect 1195 -1985 1205 -1415
rect 1115 -1995 1205 -1985
rect -95 -2415 -5 -2405
rect -95 -2985 -85 -2415
rect -65 -2985 -35 -2415
rect -15 -2985 -5 -2415
rect -95 -2995 -5 -2985
rect 55 -2415 95 -2405
rect 55 -2985 65 -2415
rect 85 -2985 95 -2415
rect 55 -2995 95 -2985
rect 155 -2415 195 -2405
rect 155 -2985 165 -2415
rect 185 -2985 195 -2415
rect 155 -2995 195 -2985
rect 255 -2415 295 -2405
rect 255 -2985 265 -2415
rect 285 -2985 295 -2415
rect 255 -2995 295 -2985
rect 355 -2415 395 -2405
rect 355 -2985 365 -2415
rect 385 -2985 395 -2415
rect 355 -2995 395 -2985
rect 435 -2415 475 -2405
rect 435 -2985 445 -2415
rect 465 -2985 475 -2415
rect 435 -2995 475 -2985
rect 535 -2415 575 -2405
rect 535 -2985 545 -2415
rect 565 -2985 575 -2415
rect 535 -2995 575 -2985
rect 635 -2415 675 -2405
rect 635 -2985 645 -2415
rect 665 -2985 675 -2415
rect 635 -2995 675 -2985
rect 715 -2415 755 -2405
rect 715 -2985 725 -2415
rect 745 -2985 755 -2415
rect 715 -2995 755 -2985
rect 815 -2415 855 -2405
rect 815 -2985 825 -2415
rect 845 -2985 855 -2415
rect 815 -2995 855 -2985
rect 915 -2415 955 -2405
rect 915 -2985 925 -2415
rect 945 -2985 955 -2415
rect 915 -2995 955 -2985
rect 1015 -2415 1055 -2405
rect 1015 -2985 1025 -2415
rect 1045 -2985 1055 -2415
rect 1015 -2995 1055 -2985
rect 1115 -2415 1205 -2405
rect 1115 -2985 1125 -2415
rect 1145 -2985 1175 -2415
rect 1195 -2985 1205 -2415
rect 1115 -2995 1205 -2985
<< end >>
