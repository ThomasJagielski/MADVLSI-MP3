magic
tech sky130A
timestamp 1615822302
<< nwell >>
rect -220 -935 1330 635
<< nmos >>
rect -100 -1750 -50 -1150
rect 0 -1750 50 -1150
rect 100 -1750 150 -1150
rect 200 -1750 250 -1150
rect 300 -1750 350 -1150
rect 480 -1750 530 -1150
rect 580 -1750 630 -1150
rect 760 -1750 810 -1150
rect 860 -1750 910 -1150
rect 960 -1750 1010 -1150
rect 1060 -1750 1110 -1150
rect 1160 -1750 1210 -1150
rect -100 -2575 -50 -1975
rect 0 -2575 50 -1975
rect 100 -2575 150 -1975
rect 200 -2575 250 -1975
rect 300 -2575 350 -1975
rect 480 -2575 530 -1975
rect 580 -2575 630 -1975
rect 760 -2575 810 -1975
rect 860 -2575 910 -1975
rect 960 -2575 1010 -1975
rect 1060 -2575 1110 -1975
rect 1160 -2575 1210 -1975
<< pmos >>
rect -100 15 -50 615
rect 0 15 50 615
rect 100 15 150 615
rect 280 15 330 615
rect 380 15 430 615
rect 480 15 530 615
rect 580 15 630 615
rect 680 15 730 615
rect 780 15 830 615
rect 960 15 1010 615
rect 1060 15 1110 615
rect 1160 15 1210 615
rect -100 -915 -50 -315
rect 0 -915 50 -315
rect 100 -915 150 -315
rect 200 -915 250 -315
rect 300 -915 350 -315
rect 480 -915 530 -315
rect 580 -915 630 -315
rect 760 -915 810 -315
rect 860 -915 910 -315
rect 960 -915 1010 -315
rect 1060 -915 1110 -315
rect 1160 -915 1210 -315
<< ndiff >>
rect -150 -1165 -100 -1150
rect -150 -1735 -135 -1165
rect -115 -1735 -100 -1165
rect -150 -1750 -100 -1735
rect -50 -1165 0 -1150
rect -50 -1735 -35 -1165
rect -15 -1735 0 -1165
rect -50 -1750 0 -1735
rect 50 -1165 100 -1150
rect 50 -1735 65 -1165
rect 85 -1735 100 -1165
rect 50 -1750 100 -1735
rect 150 -1165 200 -1150
rect 150 -1735 165 -1165
rect 185 -1735 200 -1165
rect 150 -1750 200 -1735
rect 250 -1165 300 -1150
rect 250 -1735 265 -1165
rect 285 -1735 300 -1165
rect 250 -1750 300 -1735
rect 350 -1165 400 -1150
rect 350 -1735 365 -1165
rect 385 -1735 400 -1165
rect 350 -1750 400 -1735
rect 430 -1165 480 -1150
rect 430 -1735 445 -1165
rect 465 -1735 480 -1165
rect 430 -1750 480 -1735
rect 530 -1165 580 -1150
rect 530 -1735 545 -1165
rect 565 -1735 580 -1165
rect 530 -1750 580 -1735
rect 630 -1165 680 -1150
rect 630 -1735 645 -1165
rect 665 -1735 680 -1165
rect 630 -1750 680 -1735
rect 710 -1165 760 -1150
rect 710 -1735 725 -1165
rect 745 -1735 760 -1165
rect 710 -1750 760 -1735
rect 810 -1165 860 -1150
rect 810 -1735 825 -1165
rect 845 -1735 860 -1165
rect 810 -1750 860 -1735
rect 910 -1165 960 -1150
rect 910 -1735 925 -1165
rect 945 -1735 960 -1165
rect 910 -1750 960 -1735
rect 1010 -1165 1060 -1150
rect 1010 -1735 1025 -1165
rect 1045 -1735 1060 -1165
rect 1010 -1750 1060 -1735
rect 1110 -1165 1160 -1150
rect 1110 -1735 1125 -1165
rect 1145 -1735 1160 -1165
rect 1110 -1750 1160 -1735
rect 1210 -1165 1260 -1150
rect 1210 -1735 1225 -1165
rect 1245 -1735 1260 -1165
rect 1210 -1750 1260 -1735
rect -150 -1990 -100 -1975
rect -150 -2560 -135 -1990
rect -115 -2560 -100 -1990
rect -150 -2575 -100 -2560
rect -50 -1990 0 -1975
rect -50 -2560 -35 -1990
rect -15 -2560 0 -1990
rect -50 -2575 0 -2560
rect 50 -1990 100 -1975
rect 50 -2560 65 -1990
rect 85 -2560 100 -1990
rect 50 -2575 100 -2560
rect 150 -1990 200 -1975
rect 150 -2560 165 -1990
rect 185 -2560 200 -1990
rect 150 -2575 200 -2560
rect 250 -1990 300 -1975
rect 250 -2560 265 -1990
rect 285 -2560 300 -1990
rect 250 -2575 300 -2560
rect 350 -1990 400 -1975
rect 350 -2560 365 -1990
rect 385 -2560 400 -1990
rect 350 -2575 400 -2560
rect 430 -1990 480 -1975
rect 430 -2560 445 -1990
rect 465 -2560 480 -1990
rect 430 -2575 480 -2560
rect 530 -1990 580 -1975
rect 530 -2560 545 -1990
rect 565 -2560 580 -1990
rect 530 -2575 580 -2560
rect 630 -1990 680 -1975
rect 630 -2560 645 -1990
rect 665 -2560 680 -1990
rect 630 -2575 680 -2560
rect 710 -1990 760 -1975
rect 710 -2560 725 -1990
rect 745 -2560 760 -1990
rect 710 -2575 760 -2560
rect 810 -1990 860 -1975
rect 810 -2560 825 -1990
rect 845 -2560 860 -1990
rect 810 -2575 860 -2560
rect 910 -1990 960 -1975
rect 910 -2560 925 -1990
rect 945 -2560 960 -1990
rect 910 -2575 960 -2560
rect 1010 -1990 1060 -1975
rect 1010 -2560 1025 -1990
rect 1045 -2560 1060 -1990
rect 1010 -2575 1060 -2560
rect 1110 -1990 1160 -1975
rect 1110 -2560 1125 -1990
rect 1145 -2560 1160 -1990
rect 1110 -2575 1160 -2560
rect 1210 -1990 1260 -1975
rect 1210 -2560 1225 -1990
rect 1245 -2560 1260 -1990
rect 1210 -2575 1260 -2560
<< pdiff >>
rect -150 600 -100 615
rect -150 30 -135 600
rect -115 30 -100 600
rect -150 15 -100 30
rect -50 600 0 615
rect -50 30 -35 600
rect -15 30 0 600
rect -50 15 0 30
rect 50 600 100 615
rect 50 30 65 600
rect 85 30 100 600
rect 50 15 100 30
rect 150 600 200 615
rect 150 30 165 600
rect 185 30 200 600
rect 150 15 200 30
rect 230 600 280 615
rect 230 30 245 600
rect 265 30 280 600
rect 230 15 280 30
rect 330 600 380 615
rect 330 30 345 600
rect 365 30 380 600
rect 330 15 380 30
rect 430 600 480 615
rect 430 30 445 600
rect 465 30 480 600
rect 430 15 480 30
rect 530 600 580 615
rect 530 30 545 600
rect 565 30 580 600
rect 530 15 580 30
rect 630 600 680 615
rect 630 30 645 600
rect 665 30 680 600
rect 630 15 680 30
rect 730 600 780 615
rect 730 30 745 600
rect 765 30 780 600
rect 730 15 780 30
rect 830 600 880 615
rect 830 30 845 600
rect 865 30 880 600
rect 830 15 880 30
rect 910 600 960 615
rect 910 30 925 600
rect 945 30 960 600
rect 910 15 960 30
rect 1010 600 1060 615
rect 1010 30 1025 600
rect 1045 30 1060 600
rect 1010 15 1060 30
rect 1110 600 1160 615
rect 1110 30 1125 600
rect 1145 30 1160 600
rect 1110 15 1160 30
rect 1210 600 1260 615
rect 1210 30 1225 600
rect 1245 30 1260 600
rect 1210 15 1260 30
rect -150 -330 -100 -315
rect -150 -900 -135 -330
rect -115 -900 -100 -330
rect -150 -915 -100 -900
rect -50 -330 0 -315
rect -50 -900 -35 -330
rect -15 -900 0 -330
rect -50 -915 0 -900
rect 50 -330 100 -315
rect 50 -900 65 -330
rect 85 -900 100 -330
rect 50 -915 100 -900
rect 150 -330 200 -315
rect 150 -900 165 -330
rect 185 -900 200 -330
rect 150 -915 200 -900
rect 250 -330 300 -315
rect 250 -900 265 -330
rect 285 -900 300 -330
rect 250 -915 300 -900
rect 350 -330 400 -315
rect 350 -900 365 -330
rect 385 -900 400 -330
rect 350 -915 400 -900
rect 430 -330 480 -315
rect 430 -900 445 -330
rect 465 -900 480 -330
rect 430 -915 480 -900
rect 530 -330 580 -315
rect 530 -900 545 -330
rect 565 -900 580 -330
rect 530 -915 580 -900
rect 630 -330 680 -315
rect 630 -900 645 -330
rect 665 -900 680 -330
rect 630 -915 680 -900
rect 710 -330 760 -315
rect 710 -900 725 -330
rect 745 -900 760 -330
rect 710 -915 760 -900
rect 810 -330 860 -315
rect 810 -900 825 -330
rect 845 -900 860 -330
rect 810 -915 860 -900
rect 910 -330 960 -315
rect 910 -900 925 -330
rect 945 -900 960 -330
rect 910 -915 960 -900
rect 1010 -330 1060 -315
rect 1010 -900 1025 -330
rect 1045 -900 1060 -330
rect 1010 -915 1060 -900
rect 1110 -330 1160 -315
rect 1110 -900 1125 -330
rect 1145 -900 1160 -330
rect 1110 -915 1160 -900
rect 1210 -330 1260 -315
rect 1210 -900 1225 -330
rect 1245 -900 1260 -330
rect 1210 -915 1260 -900
<< ndiffc >>
rect -135 -1735 -115 -1165
rect -35 -1735 -15 -1165
rect 65 -1735 85 -1165
rect 165 -1735 185 -1165
rect 265 -1735 285 -1165
rect 365 -1735 385 -1165
rect 445 -1735 465 -1165
rect 545 -1735 565 -1165
rect 645 -1735 665 -1165
rect 725 -1735 745 -1165
rect 825 -1735 845 -1165
rect 925 -1735 945 -1165
rect 1025 -1735 1045 -1165
rect 1125 -1735 1145 -1165
rect 1225 -1735 1245 -1165
rect -135 -2560 -115 -1990
rect -35 -2560 -15 -1990
rect 65 -2560 85 -1990
rect 165 -2560 185 -1990
rect 265 -2560 285 -1990
rect 365 -2560 385 -1990
rect 445 -2560 465 -1990
rect 545 -2560 565 -1990
rect 645 -2560 665 -1990
rect 725 -2560 745 -1990
rect 825 -2560 845 -1990
rect 925 -2560 945 -1990
rect 1025 -2560 1045 -1990
rect 1125 -2560 1145 -1990
rect 1225 -2560 1245 -1990
<< pdiffc >>
rect -135 30 -115 600
rect -35 30 -15 600
rect 65 30 85 600
rect 165 30 185 600
rect 245 30 265 600
rect 345 30 365 600
rect 445 30 465 600
rect 545 30 565 600
rect 645 30 665 600
rect 745 30 765 600
rect 845 30 865 600
rect 925 30 945 600
rect 1025 30 1045 600
rect 1125 30 1145 600
rect 1225 30 1245 600
rect -135 -900 -115 -330
rect -35 -900 -15 -330
rect 65 -900 85 -330
rect 165 -900 185 -330
rect 265 -900 285 -330
rect 365 -900 385 -330
rect 445 -900 465 -330
rect 545 -900 565 -330
rect 645 -900 665 -330
rect 725 -900 745 -330
rect 825 -900 845 -330
rect 925 -900 945 -330
rect 1025 -900 1045 -330
rect 1125 -900 1145 -330
rect 1225 -900 1245 -330
<< psubdiff >>
rect -200 -1165 -150 -1150
rect -200 -1735 -185 -1165
rect -165 -1735 -150 -1165
rect -200 -1750 -150 -1735
rect 1260 -1165 1310 -1150
rect 1260 -1735 1275 -1165
rect 1295 -1735 1310 -1165
rect 1260 -1750 1310 -1735
rect -200 -1990 -150 -1975
rect -200 -2560 -185 -1990
rect -165 -2560 -150 -1990
rect -200 -2575 -150 -2560
rect 1260 -1990 1310 -1975
rect 1260 -2560 1275 -1990
rect 1295 -2560 1310 -1990
rect 1260 -2575 1310 -2560
<< nsubdiff >>
rect -200 600 -150 615
rect -200 30 -185 600
rect -165 30 -150 600
rect -200 15 -150 30
rect 1260 600 1310 615
rect 1260 30 1275 600
rect 1295 30 1310 600
rect 1260 15 1310 30
rect -200 -330 -150 -315
rect -200 -900 -185 -330
rect -165 -900 -150 -330
rect -200 -915 -150 -900
rect 1260 -330 1310 -315
rect 1260 -900 1275 -330
rect 1295 -900 1310 -330
rect 1260 -915 1310 -900
<< psubdiffcont >>
rect -185 -1735 -165 -1165
rect 1275 -1735 1295 -1165
rect -185 -2560 -165 -1990
rect 1275 -2560 1295 -1990
<< nsubdiffcont >>
rect -185 30 -165 600
rect 1275 30 1295 600
rect -185 -900 -165 -330
rect 1275 -900 1295 -330
<< poly >>
rect 1060 660 1110 670
rect 1060 640 1080 660
rect 1100 640 1110 660
rect -100 615 -50 630
rect 0 615 50 630
rect 100 615 150 630
rect 280 615 330 630
rect 380 615 430 630
rect 480 615 530 630
rect 580 615 630 630
rect 680 615 730 630
rect 780 615 830 630
rect 960 615 1010 630
rect 1060 615 1110 640
rect 1160 615 1210 630
rect -100 0 -50 15
rect -150 -10 -50 0
rect -150 -30 -140 -10
rect -120 -30 -50 -10
rect -150 -40 -50 -30
rect 0 5 50 15
rect 100 5 150 15
rect 280 5 330 15
rect 380 5 430 15
rect 480 5 530 15
rect 580 5 630 15
rect 680 5 730 15
rect 780 5 830 15
rect 960 5 1010 15
rect 1060 5 1110 15
rect 0 -10 1110 5
rect 1160 0 1210 15
rect 0 -65 15 -10
rect 1160 -15 1260 0
rect 1160 -35 1230 -15
rect 1250 -35 1260 -15
rect 1160 -45 1260 -35
rect -150 -75 15 -65
rect -150 -95 -140 -75
rect -120 -80 15 -75
rect -120 -95 -110 -80
rect -150 -105 -110 -95
rect -45 -270 -5 -260
rect -45 -290 -35 -270
rect -15 -290 -5 -270
rect 255 -270 295 -260
rect 255 -285 265 -270
rect 100 -290 265 -285
rect 285 -285 295 -270
rect 535 -270 575 -260
rect 285 -290 350 -285
rect 535 -290 545 -270
rect 565 -290 575 -270
rect 815 -270 855 -260
rect 815 -285 825 -270
rect 760 -290 825 -285
rect 845 -285 855 -270
rect 1115 -270 1155 -260
rect 845 -290 1010 -285
rect 1115 -290 1125 -270
rect 1145 -290 1155 -270
rect -100 -305 50 -290
rect -100 -315 -50 -305
rect 0 -315 50 -305
rect 100 -300 350 -290
rect 100 -315 150 -300
rect 200 -315 250 -300
rect 300 -315 350 -300
rect 480 -305 630 -290
rect 480 -315 530 -305
rect 580 -315 630 -305
rect 760 -300 1010 -290
rect 760 -315 810 -300
rect 860 -315 910 -300
rect 960 -315 1010 -300
rect 1060 -305 1210 -290
rect 1060 -315 1110 -305
rect 1160 -315 1210 -305
rect -100 -930 -50 -915
rect 0 -930 50 -915
rect 100 -1045 150 -915
rect 200 -930 250 -915
rect 300 -930 350 -915
rect 480 -930 530 -915
rect 580 -980 630 -915
rect 760 -930 810 -915
rect 860 -930 910 -915
rect 960 -930 1010 -915
rect 1060 -930 1110 -915
rect 1160 -930 1210 -915
rect 580 -1000 595 -980
rect 615 -1000 630 -980
rect 580 -1010 630 -1000
rect 100 -1065 115 -1045
rect 135 -1065 150 -1045
rect 100 -1075 150 -1065
rect 475 -1045 515 -1035
rect 475 -1065 485 -1045
rect 505 -1060 515 -1045
rect 595 -1045 635 -1035
rect 595 -1060 605 -1045
rect 505 -1065 605 -1060
rect 625 -1065 635 -1045
rect 1115 -1040 1155 -1030
rect 1115 -1055 1125 -1040
rect 475 -1075 635 -1065
rect 995 -1060 1125 -1055
rect 1145 -1060 1155 -1040
rect 995 -1070 1155 -1060
rect -45 -1105 -5 -1095
rect -45 -1120 -35 -1105
rect -100 -1125 -35 -1120
rect -15 -1120 -5 -1105
rect 355 -1105 395 -1095
rect 355 -1120 365 -1105
rect -15 -1125 50 -1120
rect -100 -1135 50 -1125
rect -100 -1150 -50 -1135
rect 0 -1150 50 -1135
rect 100 -1125 365 -1120
rect 385 -1120 395 -1105
rect 715 -1105 755 -1095
rect 715 -1120 725 -1105
rect 385 -1125 725 -1120
rect 745 -1120 755 -1105
rect 995 -1120 1010 -1070
rect 1115 -1105 1155 -1095
rect 1115 -1120 1125 -1105
rect 745 -1125 1010 -1120
rect 100 -1135 1010 -1125
rect 100 -1150 150 -1135
rect 200 -1150 250 -1135
rect 300 -1150 350 -1135
rect 480 -1150 530 -1135
rect 580 -1150 630 -1135
rect 760 -1150 810 -1135
rect 860 -1150 910 -1135
rect 960 -1150 1010 -1135
rect 1060 -1125 1125 -1120
rect 1145 -1120 1155 -1105
rect 1145 -1125 1210 -1120
rect 1060 -1135 1210 -1125
rect 1060 -1150 1110 -1135
rect 1160 -1150 1210 -1135
rect -100 -1765 -50 -1750
rect 0 -1765 50 -1750
rect 100 -1765 150 -1750
rect 200 -1765 250 -1750
rect 300 -1765 350 -1750
rect 480 -1765 530 -1750
rect 580 -1765 630 -1750
rect 760 -1765 810 -1750
rect 860 -1765 910 -1750
rect 960 -1765 1010 -1750
rect 1060 -1765 1110 -1750
rect 1160 -1765 1210 -1750
rect 235 -1920 295 -1910
rect -45 -1930 -5 -1920
rect -45 -1945 -35 -1930
rect -100 -1950 -35 -1945
rect -15 -1945 -5 -1930
rect 235 -1940 265 -1920
rect 285 -1930 855 -1920
rect 285 -1935 825 -1930
rect 285 -1940 350 -1935
rect 235 -1945 350 -1940
rect -15 -1950 50 -1945
rect -100 -1960 50 -1950
rect -100 -1975 -50 -1960
rect 0 -1975 50 -1960
rect 100 -1950 350 -1945
rect 100 -1960 250 -1950
rect 100 -1975 150 -1960
rect 200 -1975 250 -1960
rect 300 -1975 350 -1950
rect 760 -1950 825 -1935
rect 845 -1945 855 -1930
rect 1115 -1930 1155 -1920
rect 1115 -1945 1125 -1930
rect 845 -1950 1010 -1945
rect 760 -1960 1010 -1950
rect 480 -1975 530 -1960
rect 580 -1975 630 -1960
rect 760 -1975 810 -1960
rect 860 -1975 910 -1960
rect 960 -1975 1010 -1960
rect 1060 -1950 1125 -1945
rect 1145 -1945 1155 -1930
rect 1145 -1950 1210 -1945
rect 1060 -1960 1210 -1950
rect 1060 -1975 1110 -1960
rect 1160 -1975 1210 -1960
rect -100 -2590 -50 -2575
rect 0 -2590 50 -2575
rect 100 -2590 150 -2575
rect 200 -2590 250 -2575
rect 300 -2590 350 -2575
rect 480 -2590 530 -2575
rect 580 -2590 630 -2575
rect 760 -2590 810 -2575
rect 860 -2590 910 -2575
rect 960 -2590 1010 -2575
rect 1060 -2590 1110 -2575
rect 1160 -2590 1210 -2575
rect 480 -2600 630 -2590
rect 480 -2610 545 -2600
rect 535 -2620 545 -2610
rect 565 -2610 630 -2600
rect 565 -2620 575 -2610
rect 535 -2630 575 -2620
<< polycont >>
rect 1080 640 1100 660
rect -140 -30 -120 -10
rect 1230 -35 1250 -15
rect -140 -95 -120 -75
rect -35 -290 -15 -270
rect 265 -290 285 -270
rect 545 -290 565 -270
rect 825 -290 845 -270
rect 1125 -290 1145 -270
rect 595 -1000 615 -980
rect 115 -1065 135 -1045
rect 485 -1065 505 -1045
rect 605 -1065 625 -1045
rect 1125 -1060 1145 -1040
rect -35 -1125 -15 -1105
rect 365 -1125 385 -1105
rect 725 -1125 745 -1105
rect 1125 -1125 1145 -1105
rect -35 -1950 -15 -1930
rect 265 -1940 285 -1920
rect 825 -1950 845 -1930
rect 1125 -1950 1145 -1930
rect 545 -2620 565 -2600
<< locali >>
rect 1060 660 1310 670
rect 1060 640 1080 660
rect 1100 640 1310 660
rect 1060 630 1310 640
rect -195 600 -105 610
rect -195 30 -185 600
rect -165 30 -135 600
rect -115 30 -105 600
rect -195 20 -105 30
rect -150 -10 -105 20
rect -150 -30 -140 -10
rect -120 -30 -105 -10
rect -150 -40 -105 -30
rect -45 600 -5 610
rect -45 30 -35 600
rect -15 30 -5 600
rect -45 -65 -5 30
rect 55 600 95 610
rect 55 30 65 600
rect 85 30 95 600
rect 55 20 95 30
rect 155 600 195 610
rect 155 30 165 600
rect 185 30 195 600
rect -200 -75 -5 -65
rect -200 -95 -140 -75
rect -120 -85 -5 -75
rect -120 -95 -110 -85
rect -200 -105 -110 -95
rect 155 -125 195 30
rect 235 600 275 610
rect 235 30 245 600
rect 265 30 275 600
rect 235 -95 275 30
rect 335 600 375 610
rect 335 30 345 600
rect 365 30 375 600
rect 335 25 375 30
rect 435 600 475 610
rect 435 30 445 600
rect 465 30 475 600
rect 435 20 475 30
rect 535 600 575 610
rect 535 30 545 600
rect 565 30 575 600
rect 535 -45 575 30
rect 635 600 675 610
rect 635 30 645 600
rect 665 30 675 600
rect 635 20 675 30
rect 735 600 775 610
rect 735 30 745 600
rect 765 30 775 600
rect 735 25 775 30
rect 835 600 875 610
rect 835 30 845 600
rect 865 30 875 600
rect 535 -65 545 -45
rect 565 -65 575 -45
rect 535 -75 575 -65
rect 835 -85 875 30
rect 835 -95 845 -85
rect 235 -105 845 -95
rect 865 -105 875 -85
rect 235 -115 875 -105
rect 915 600 955 610
rect 915 30 925 600
rect 945 30 955 600
rect 155 -145 165 -125
rect 185 -135 195 -125
rect 915 -135 955 30
rect 1015 600 1055 610
rect 1015 30 1025 600
rect 1045 30 1055 600
rect 1015 20 1055 30
rect 1115 600 1155 630
rect 1115 30 1125 600
rect 1145 30 1155 600
rect 1115 20 1155 30
rect 1215 600 1305 610
rect 1215 30 1225 600
rect 1245 30 1275 600
rect 1295 30 1305 600
rect 1215 20 1305 30
rect 1215 -15 1260 20
rect 1215 -35 1230 -15
rect 1250 -35 1260 -15
rect 1215 -45 1260 -35
rect 185 -145 955 -135
rect 155 -155 955 -145
rect 255 -240 855 -220
rect -150 -270 -5 -260
rect -150 -280 -35 -270
rect -150 -320 -105 -280
rect -195 -330 -105 -320
rect -195 -900 -185 -330
rect -165 -900 -135 -330
rect -115 -900 -105 -330
rect -195 -910 -105 -900
rect -45 -290 -35 -280
rect -15 -290 -5 -270
rect -45 -330 -5 -290
rect 255 -270 395 -240
rect 255 -290 265 -270
rect 285 -290 395 -270
rect 255 -300 395 -290
rect -45 -900 -35 -330
rect -15 -900 -5 -330
rect -45 -910 -5 -900
rect 55 -330 95 -320
rect 55 -900 65 -330
rect 85 -900 95 -330
rect 55 -910 95 -900
rect 155 -330 195 -320
rect 155 -900 165 -330
rect 185 -900 195 -330
rect 155 -930 195 -900
rect 255 -330 295 -300
rect 255 -900 265 -330
rect 285 -900 295 -330
rect 255 -910 295 -900
rect 355 -330 395 -300
rect 535 -270 575 -260
rect 535 -290 545 -270
rect 565 -290 575 -270
rect 355 -900 365 -330
rect 385 -900 395 -330
rect 355 -910 395 -900
rect 435 -330 475 -320
rect 435 -900 445 -330
rect 465 -900 475 -330
rect 435 -930 475 -900
rect 535 -330 575 -290
rect 715 -270 855 -240
rect 715 -290 825 -270
rect 845 -290 855 -270
rect 715 -300 855 -290
rect 535 -900 545 -330
rect 565 -900 575 -330
rect 535 -910 575 -900
rect 635 -330 675 -320
rect 635 -900 645 -330
rect 665 -900 675 -330
rect 635 -930 675 -900
rect 715 -330 755 -300
rect 715 -900 725 -330
rect 745 -900 755 -330
rect 715 -910 755 -900
rect 815 -330 855 -300
rect 1115 -270 1260 -260
rect 1115 -290 1125 -270
rect 1145 -280 1260 -270
rect 1145 -290 1155 -280
rect 815 -900 825 -330
rect 845 -900 855 -330
rect 815 -910 855 -900
rect 915 -330 955 -320
rect 915 -900 925 -330
rect 945 -900 955 -330
rect 915 -930 955 -900
rect 1015 -330 1055 -320
rect 1015 -900 1025 -330
rect 1045 -900 1055 -330
rect 1015 -910 1055 -900
rect 1115 -330 1155 -290
rect 1115 -900 1125 -330
rect 1145 -900 1155 -330
rect 1115 -910 1155 -900
rect 1215 -320 1260 -280
rect 1215 -330 1305 -320
rect 1215 -900 1225 -330
rect 1245 -900 1275 -330
rect 1295 -900 1305 -330
rect 1215 -910 1305 -900
rect 155 -950 955 -930
rect 535 -980 1310 -970
rect 535 -1000 595 -980
rect 615 -990 1310 -980
rect 615 -1000 630 -990
rect 535 -1010 630 -1000
rect 100 -1045 150 -1035
rect 100 -1055 115 -1045
rect 55 -1065 115 -1055
rect 135 -1055 150 -1045
rect 475 -1045 515 -1035
rect 475 -1055 485 -1045
rect 135 -1065 485 -1055
rect 505 -1065 515 -1045
rect 55 -1075 515 -1065
rect -150 -1105 -5 -1095
rect -150 -1115 -35 -1105
rect -150 -1155 -105 -1115
rect -195 -1165 -105 -1155
rect -195 -1735 -185 -1165
rect -165 -1735 -135 -1165
rect -115 -1735 -105 -1165
rect -195 -1745 -105 -1735
rect -45 -1125 -35 -1115
rect -15 -1125 -5 -1105
rect -45 -1165 -5 -1125
rect -45 -1735 -35 -1165
rect -15 -1735 -5 -1165
rect -45 -1745 -5 -1735
rect 55 -1165 95 -1075
rect 355 -1105 395 -1095
rect 355 -1125 365 -1105
rect 385 -1125 395 -1105
rect 55 -1735 65 -1165
rect 85 -1735 95 -1165
rect 55 -1745 95 -1735
rect 155 -1165 195 -1155
rect 155 -1735 165 -1165
rect 185 -1735 195 -1165
rect 155 -1745 195 -1735
rect 255 -1165 295 -1155
rect 255 -1735 265 -1165
rect 285 -1735 295 -1165
rect 255 -1830 295 -1735
rect 355 -1165 395 -1125
rect 355 -1735 365 -1165
rect 385 -1735 395 -1165
rect 355 -1745 395 -1735
rect 435 -1165 475 -1155
rect 435 -1735 445 -1165
rect 465 -1735 475 -1165
rect 435 -1830 475 -1735
rect 535 -1165 575 -1010
rect 595 -1045 635 -1035
rect 595 -1065 605 -1045
rect 625 -1055 635 -1045
rect 1115 -1040 1155 -1030
rect 625 -1065 1055 -1055
rect 595 -1075 1055 -1065
rect 1115 -1060 1125 -1040
rect 1145 -1050 1155 -1040
rect 1145 -1060 1310 -1050
rect 1115 -1070 1310 -1060
rect 715 -1105 755 -1095
rect 715 -1125 725 -1105
rect 745 -1125 755 -1105
rect 535 -1735 545 -1165
rect 565 -1735 575 -1165
rect 535 -1745 575 -1735
rect 635 -1165 675 -1155
rect 635 -1735 645 -1165
rect 665 -1735 675 -1165
rect 635 -1830 675 -1735
rect 715 -1165 755 -1125
rect 715 -1735 725 -1165
rect 745 -1735 755 -1165
rect 715 -1745 755 -1735
rect 815 -1165 855 -1155
rect 815 -1735 825 -1165
rect 845 -1735 855 -1165
rect 815 -1745 855 -1735
rect 915 -1165 955 -1155
rect 915 -1735 925 -1165
rect 945 -1735 955 -1165
rect 915 -1745 955 -1735
rect 1015 -1165 1055 -1075
rect 1015 -1735 1025 -1165
rect 1045 -1735 1055 -1165
rect 1015 -1745 1055 -1735
rect 1115 -1105 1260 -1095
rect 1115 -1125 1125 -1105
rect 1145 -1115 1260 -1105
rect 1145 -1125 1155 -1115
rect 1115 -1165 1155 -1125
rect 1115 -1735 1125 -1165
rect 1145 -1735 1155 -1165
rect 1115 -1745 1155 -1735
rect 1215 -1155 1260 -1115
rect 1215 -1165 1305 -1155
rect 1215 -1735 1225 -1165
rect 1245 -1735 1275 -1165
rect 1295 -1735 1305 -1165
rect 1215 -1745 1305 -1735
rect 810 -1830 855 -1745
rect 255 -1850 855 -1830
rect 155 -1890 955 -1870
rect -150 -1930 -5 -1920
rect -150 -1940 -35 -1930
rect -150 -1980 -105 -1940
rect -45 -1950 -35 -1940
rect -15 -1950 -5 -1930
rect -45 -1960 -5 -1950
rect -195 -1990 -105 -1980
rect -195 -2560 -185 -1990
rect -165 -2560 -135 -1990
rect -115 -2560 -105 -1990
rect -195 -2570 -105 -2560
rect -45 -1990 -5 -1980
rect -45 -2560 -35 -1990
rect -15 -2560 -5 -1990
rect -45 -2570 -5 -2560
rect 55 -1990 95 -1980
rect 55 -2560 65 -1990
rect 85 -2560 95 -1990
rect 55 -2570 95 -2560
rect 155 -1990 195 -1890
rect 155 -2560 165 -1990
rect 185 -2560 195 -1990
rect 155 -2570 195 -2560
rect 255 -1920 395 -1910
rect 255 -1940 265 -1920
rect 285 -1940 395 -1920
rect 255 -1950 395 -1940
rect 255 -1990 295 -1950
rect 255 -2560 265 -1990
rect 285 -2560 295 -1990
rect 255 -2570 295 -2560
rect 355 -1990 395 -1950
rect 355 -2560 365 -1990
rect 385 -2560 395 -1990
rect 355 -2570 395 -2560
rect 435 -1990 475 -1890
rect 435 -2560 445 -1990
rect 465 -2560 475 -1990
rect 435 -2570 475 -2560
rect 535 -1920 575 -1910
rect 535 -1940 545 -1920
rect 565 -1940 575 -1920
rect 535 -1990 575 -1940
rect 535 -2560 545 -1990
rect 565 -2560 575 -1990
rect 535 -2600 575 -2560
rect 635 -1990 675 -1890
rect 635 -2560 645 -1990
rect 665 -2560 675 -1990
rect 635 -2570 675 -2560
rect 715 -1930 855 -1920
rect 715 -1950 825 -1930
rect 845 -1950 855 -1930
rect 715 -1960 855 -1950
rect 715 -1990 755 -1960
rect 715 -2560 725 -1990
rect 745 -2560 755 -1990
rect 715 -2570 755 -2560
rect 815 -1990 855 -1960
rect 815 -2560 825 -1990
rect 845 -2560 855 -1990
rect 815 -2570 855 -2560
rect 915 -1990 955 -1890
rect 1115 -1930 1260 -1920
rect 1115 -1950 1125 -1930
rect 1145 -1945 1260 -1930
rect 1145 -1950 1155 -1945
rect 915 -2560 925 -1990
rect 945 -2560 955 -1990
rect 915 -2570 955 -2560
rect 1015 -1990 1055 -1980
rect 1015 -2560 1025 -1990
rect 1045 -2560 1055 -1990
rect 1015 -2570 1055 -2560
rect 1115 -1990 1155 -1950
rect 1115 -2560 1125 -1990
rect 1145 -2560 1155 -1990
rect 1115 -2570 1155 -2560
rect 1215 -1980 1260 -1945
rect 1215 -1990 1305 -1980
rect 1215 -2560 1225 -1990
rect 1245 -2560 1275 -1990
rect 1295 -2560 1305 -1990
rect 1215 -2570 1305 -2560
rect 535 -2620 545 -2600
rect 565 -2610 575 -2600
rect 565 -2620 1310 -2610
rect 535 -2630 1310 -2620
<< viali >>
rect -185 30 -165 600
rect -135 30 -115 600
rect 65 30 85 600
rect 345 30 365 600
rect 745 30 765 600
rect 545 -65 565 -45
rect 845 -105 865 -85
rect 165 -145 185 -125
rect 1025 30 1045 600
rect 1225 30 1245 600
rect 1275 30 1295 600
rect -185 -900 -165 -330
rect -135 -900 -115 -330
rect -35 -900 -15 -330
rect 65 -900 85 -330
rect 1025 -900 1045 -330
rect 1125 -900 1145 -330
rect 1225 -900 1245 -330
rect 1275 -900 1295 -330
rect -185 -1735 -165 -1165
rect -135 -1735 -115 -1165
rect -35 -1735 -15 -1165
rect 365 -1125 385 -1105
rect 265 -1735 285 -1165
rect 825 -1735 845 -1165
rect 1125 -1735 1145 -1165
rect 1225 -1735 1245 -1165
rect 1275 -1735 1295 -1165
rect -185 -2560 -165 -1990
rect -135 -2560 -115 -1990
rect -35 -2560 -15 -1990
rect 65 -2560 85 -1990
rect 265 -1940 285 -1920
rect 545 -1940 565 -1920
rect 1025 -2560 1045 -1990
rect 1125 -2560 1145 -1990
rect 1225 -2560 1245 -1990
rect 1275 -2560 1295 -1990
<< metal1 >>
rect -200 600 1310 610
rect -200 30 -185 600
rect -165 30 -135 600
rect -115 30 65 600
rect 85 30 345 600
rect 365 30 745 600
rect 765 30 1025 600
rect 1045 30 1225 600
rect 1245 30 1275 600
rect 1295 30 1310 600
rect -200 20 1310 30
rect -200 -330 95 20
rect 535 -45 575 -35
rect 535 -65 545 -45
rect 565 -65 575 -45
rect -200 -900 -185 -330
rect -165 -900 -135 -330
rect -115 -900 -35 -330
rect -15 -900 65 -330
rect 85 -900 95 -330
rect -200 -910 95 -900
rect 155 -125 195 -115
rect 155 -145 165 -125
rect 185 -145 195 -125
rect 155 -1095 195 -145
rect 155 -1105 395 -1095
rect 155 -1125 365 -1105
rect 385 -1125 395 -1105
rect 355 -1135 395 -1125
rect -200 -1165 295 -1155
rect -200 -1735 -185 -1165
rect -165 -1735 -135 -1165
rect -115 -1735 -35 -1165
rect -15 -1735 265 -1165
rect 285 -1735 295 -1165
rect -200 -1745 295 -1735
rect -200 -1980 200 -1745
rect 535 -1810 575 -65
rect 835 -85 875 -75
rect 835 -105 845 -85
rect 865 -105 875 -85
rect 835 -1005 875 -105
rect 1015 -330 1310 20
rect 1015 -900 1025 -330
rect 1045 -900 1125 -330
rect 1145 -900 1225 -330
rect 1245 -900 1275 -330
rect 1295 -900 1310 -330
rect 1015 -910 1310 -900
rect 255 -1850 575 -1810
rect 635 -1035 875 -1005
rect 255 -1920 295 -1850
rect 635 -1910 675 -1035
rect 815 -1165 1310 -1155
rect 815 -1735 825 -1165
rect 845 -1735 1125 -1165
rect 1145 -1735 1225 -1165
rect 1245 -1735 1275 -1165
rect 1295 -1735 1310 -1165
rect 815 -1745 1310 -1735
rect 255 -1940 265 -1920
rect 285 -1940 295 -1920
rect 255 -1950 295 -1940
rect 535 -1920 675 -1910
rect 535 -1940 545 -1920
rect 565 -1940 675 -1920
rect 535 -1950 675 -1940
rect 910 -1980 1310 -1745
rect -200 -1990 1310 -1980
rect -200 -2560 -185 -1990
rect -165 -2560 -135 -1990
rect -115 -2560 -35 -1990
rect -15 -2560 65 -1990
rect 85 -2560 1025 -1990
rect 1045 -2560 1125 -1990
rect 1145 -2560 1225 -1990
rect 1245 -2560 1275 -1990
rect 1295 -2560 1310 -1990
rect -200 -2570 1310 -2560
<< labels >>
rlabel locali -200 -85 -200 -85 7 Vbp
port 3 w
rlabel metal1 -200 315 -200 315 7 VP
port 1 w
rlabel metal1 -200 -2275 -200 -2275 7 VN
port 2 w
rlabel locali 1310 -2620 1310 -2620 3 Vcn
port 4 e
rlabel locali 1310 -1060 1310 -1060 3 Vbn
port 5 e
rlabel locali 1310 -980 1310 -980 3 Vcp
port 6 e
<< end >>
