magic
tech sky130A
timestamp 1615693684
<< nwell >>
rect -135 -825 1055 745
<< nmos >>
rect -15 -2465 35 -1865
rect 85 -2465 135 -1865
rect 185 -2465 235 -1865
rect 285 -2465 335 -1865
rect 385 -2465 435 -1865
rect 485 -2465 535 -1865
rect 585 -2465 635 -1865
rect 685 -2465 735 -1865
rect 785 -2465 835 -1865
rect 885 -2465 935 -1865
<< pmos >>
rect -15 575 35 725
rect 85 575 135 725
rect 185 575 235 725
rect 285 575 335 725
rect 385 575 435 725
rect 485 575 535 725
rect 585 575 635 725
rect 685 575 735 725
rect 785 575 835 725
rect 885 575 935 725
rect -15 75 35 375
rect 85 75 135 375
rect 185 75 235 375
rect 285 75 335 375
rect 385 75 435 375
rect 485 75 535 375
rect 585 75 635 375
rect 685 75 735 375
rect 785 75 835 375
rect 885 75 935 375
rect -15 -805 35 -205
rect 85 -805 135 -205
rect 185 -805 235 -205
rect 285 -805 335 -205
rect 385 -805 435 -205
rect 485 -805 535 -205
rect 585 -805 635 -205
rect 685 -805 735 -205
rect 785 -805 835 -205
rect 885 -805 935 -205
<< ndiff >>
rect -65 -1880 -15 -1865
rect -65 -2450 -50 -1880
rect -30 -2450 -15 -1880
rect -65 -2465 -15 -2450
rect 35 -1880 85 -1865
rect 35 -2450 50 -1880
rect 70 -2450 85 -1880
rect 35 -2465 85 -2450
rect 135 -1880 185 -1865
rect 135 -2450 150 -1880
rect 170 -2450 185 -1880
rect 135 -2465 185 -2450
rect 235 -1880 285 -1865
rect 235 -2450 250 -1880
rect 270 -2450 285 -1880
rect 235 -2465 285 -2450
rect 335 -1880 385 -1865
rect 335 -2450 350 -1880
rect 370 -2450 385 -1880
rect 335 -2465 385 -2450
rect 435 -1880 485 -1865
rect 435 -2450 450 -1880
rect 470 -2450 485 -1880
rect 435 -2465 485 -2450
rect 535 -1880 585 -1865
rect 535 -2450 550 -1880
rect 570 -2450 585 -1880
rect 535 -2465 585 -2450
rect 635 -1880 685 -1865
rect 635 -2450 650 -1880
rect 670 -2450 685 -1880
rect 635 -2465 685 -2450
rect 735 -1880 785 -1865
rect 735 -2450 750 -1880
rect 770 -2450 785 -1880
rect 735 -2465 785 -2450
rect 835 -1880 885 -1865
rect 835 -2450 850 -1880
rect 870 -2450 885 -1880
rect 835 -2465 885 -2450
rect 935 -1880 985 -1865
rect 935 -2450 950 -1880
rect 970 -2450 985 -1880
rect 935 -2465 985 -2450
<< pdiff >>
rect -65 715 -15 725
rect -65 590 -50 715
rect -30 590 -15 715
rect -65 575 -15 590
rect 35 715 85 725
rect 35 590 50 715
rect 70 590 85 715
rect 35 575 85 590
rect 135 715 185 725
rect 135 590 150 715
rect 170 590 185 715
rect 135 575 185 590
rect 235 715 285 725
rect 235 590 250 715
rect 270 590 285 715
rect 235 575 285 590
rect 335 715 385 725
rect 335 590 350 715
rect 370 590 385 715
rect 335 575 385 590
rect 435 715 485 725
rect 435 590 450 715
rect 470 590 485 715
rect 435 575 485 590
rect 535 715 585 725
rect 535 590 550 715
rect 570 590 585 715
rect 535 575 585 590
rect 635 715 685 725
rect 635 590 650 715
rect 670 590 685 715
rect 635 575 685 590
rect 735 715 785 725
rect 735 590 750 715
rect 770 590 785 715
rect 735 575 785 590
rect 835 715 885 725
rect 835 590 850 715
rect 870 590 885 715
rect 835 575 885 590
rect 935 715 985 725
rect 935 590 950 715
rect 970 590 985 715
rect 935 575 985 590
rect -65 360 -15 375
rect -65 90 -50 360
rect -30 90 -15 360
rect -65 75 -15 90
rect 35 360 85 375
rect 35 90 50 360
rect 70 90 85 360
rect 35 75 85 90
rect 135 360 185 375
rect 135 90 150 360
rect 170 90 185 360
rect 135 75 185 90
rect 235 360 285 375
rect 235 90 250 360
rect 270 90 285 360
rect 235 75 285 90
rect 335 360 385 375
rect 335 90 350 360
rect 370 90 385 360
rect 335 75 385 90
rect 435 360 485 375
rect 435 90 450 360
rect 470 90 485 360
rect 435 75 485 90
rect 535 360 585 375
rect 535 90 550 360
rect 570 90 585 360
rect 535 75 585 90
rect 635 360 685 375
rect 635 90 650 360
rect 670 90 685 360
rect 635 75 685 90
rect 735 360 785 375
rect 735 90 750 360
rect 770 90 785 360
rect 735 75 785 90
rect 835 360 885 375
rect 835 90 850 360
rect 870 90 885 360
rect 835 75 885 90
rect 935 360 985 375
rect 935 90 950 360
rect 970 90 985 360
rect 935 75 985 90
rect -65 -220 -15 -205
rect -65 -790 -50 -220
rect -30 -790 -15 -220
rect -65 -805 -15 -790
rect 35 -220 85 -205
rect 35 -790 50 -220
rect 70 -790 85 -220
rect 35 -805 85 -790
rect 135 -220 185 -205
rect 135 -790 150 -220
rect 170 -790 185 -220
rect 135 -805 185 -790
rect 235 -220 285 -205
rect 235 -790 250 -220
rect 270 -790 285 -220
rect 235 -805 285 -790
rect 335 -220 385 -205
rect 335 -790 350 -220
rect 370 -790 385 -220
rect 335 -805 385 -790
rect 435 -220 485 -205
rect 435 -790 450 -220
rect 470 -790 485 -220
rect 435 -805 485 -790
rect 535 -220 585 -205
rect 535 -790 550 -220
rect 570 -790 585 -220
rect 535 -805 585 -790
rect 635 -220 685 -205
rect 635 -790 650 -220
rect 670 -790 685 -220
rect 635 -805 685 -790
rect 735 -220 785 -205
rect 735 -790 750 -220
rect 770 -790 785 -220
rect 735 -805 785 -790
rect 835 -220 885 -205
rect 835 -790 850 -220
rect 870 -790 885 -220
rect 835 -805 885 -790
rect 935 -220 985 -205
rect 935 -790 950 -220
rect 970 -790 985 -220
rect 935 -805 985 -790
<< ndiffc >>
rect -50 -2450 -30 -1880
rect 50 -2450 70 -1880
rect 150 -2450 170 -1880
rect 250 -2450 270 -1880
rect 350 -2450 370 -1880
rect 450 -2450 470 -1880
rect 550 -2450 570 -1880
rect 650 -2450 670 -1880
rect 750 -2450 770 -1880
rect 850 -2450 870 -1880
rect 950 -2450 970 -1880
<< pdiffc >>
rect -50 590 -30 715
rect 50 590 70 715
rect 150 590 170 715
rect 250 590 270 715
rect 350 590 370 715
rect 450 590 470 715
rect 550 590 570 715
rect 650 590 670 715
rect 750 590 770 715
rect 850 590 870 715
rect 950 590 970 715
rect -50 90 -30 360
rect 50 90 70 360
rect 150 90 170 360
rect 250 90 270 360
rect 350 90 370 360
rect 450 90 470 360
rect 550 90 570 360
rect 650 90 670 360
rect 750 90 770 360
rect 850 90 870 360
rect 950 90 970 360
rect -50 -790 -30 -220
rect 50 -790 70 -220
rect 150 -790 170 -220
rect 250 -790 270 -220
rect 350 -790 370 -220
rect 450 -790 470 -220
rect 550 -790 570 -220
rect 650 -790 670 -220
rect 750 -790 770 -220
rect 850 -790 870 -220
rect 950 -790 970 -220
<< psubdiff >>
rect -115 -1880 -65 -1865
rect -115 -2450 -100 -1880
rect -80 -2450 -65 -1880
rect -115 -2465 -65 -2450
rect 985 -1880 1035 -1865
rect 985 -2450 1000 -1880
rect 1020 -2450 1035 -1880
rect 985 -2465 1035 -2450
<< nsubdiff >>
rect -115 715 -65 725
rect -115 590 -100 715
rect -80 590 -65 715
rect -115 575 -65 590
rect 985 715 1035 725
rect 985 590 1000 715
rect 1020 590 1035 715
rect 985 575 1035 590
rect -115 360 -65 375
rect -115 90 -100 360
rect -80 90 -65 360
rect -115 75 -65 90
rect 985 360 1035 375
rect 985 90 1000 360
rect 1020 90 1035 360
rect 985 75 1035 90
rect -115 -220 -65 -205
rect -115 -790 -100 -220
rect -80 -790 -65 -220
rect -115 -805 -65 -790
rect 985 -220 1035 -205
rect 985 -790 1000 -220
rect 1020 -790 1035 -220
rect 985 -805 1035 -790
<< psubdiffcont >>
rect -100 -2450 -80 -1880
rect 1000 -2450 1020 -1880
<< nsubdiffcont >>
rect -100 590 -80 715
rect 1000 590 1020 715
rect -100 90 -80 360
rect 1000 90 1020 360
rect -100 -790 -80 -220
rect 1000 -790 1020 -220
<< poly >>
rect 85 770 135 780
rect 85 750 95 770
rect 115 750 135 770
rect -15 725 35 740
rect 85 725 135 750
rect 185 725 235 740
rect 285 725 335 740
rect 385 725 435 740
rect 485 725 535 740
rect 585 725 635 740
rect 685 725 735 740
rect 785 725 835 740
rect 885 725 935 740
rect -15 560 35 575
rect -60 550 35 560
rect 85 565 135 575
rect 185 565 235 575
rect 285 565 335 575
rect 385 565 435 575
rect 485 565 535 575
rect 585 565 635 575
rect 685 565 735 575
rect 785 565 835 575
rect 85 550 835 565
rect 885 560 935 575
rect 885 550 980 560
rect -60 530 -50 550
rect -30 545 35 550
rect 885 545 950 550
rect -30 530 -20 545
rect -60 520 -20 530
rect 940 530 950 545
rect 970 530 980 550
rect 940 520 980 530
rect 885 475 925 485
rect 885 460 895 475
rect 820 455 895 460
rect 915 455 925 475
rect 820 445 925 455
rect 820 430 835 445
rect -60 420 -20 430
rect -60 400 -50 420
rect -30 405 -20 420
rect 85 415 835 430
rect -30 400 35 405
rect -60 390 35 400
rect -15 375 35 390
rect 85 375 135 415
rect 185 375 235 390
rect 285 375 335 390
rect 385 375 435 415
rect 485 375 535 415
rect 585 375 635 390
rect 685 375 735 390
rect 785 375 835 415
rect 940 420 980 430
rect 940 405 950 420
rect 885 400 950 405
rect 970 400 980 420
rect 885 390 980 400
rect 885 375 935 390
rect -15 60 35 75
rect 85 60 135 75
rect 185 35 235 75
rect 285 35 335 75
rect 385 60 435 75
rect 485 60 535 75
rect 585 35 635 75
rect 685 35 735 75
rect 785 60 835 75
rect 885 60 935 75
rect 185 25 925 35
rect 185 20 895 25
rect 885 5 895 20
rect 915 5 925 25
rect 885 -5 925 5
rect 240 -15 280 -5
rect 240 -35 250 -15
rect 270 -30 280 -15
rect 640 -15 680 -5
rect 640 -30 650 -15
rect 270 -35 650 -30
rect 670 -35 680 -15
rect 240 -45 680 -35
rect 85 -135 835 -120
rect -60 -160 -20 -150
rect -60 -180 -50 -160
rect -30 -175 -20 -160
rect -30 -180 35 -175
rect -60 -190 35 -180
rect -15 -205 35 -190
rect 85 -205 135 -135
rect 185 -205 235 -190
rect 285 -205 335 -190
rect 385 -205 435 -135
rect 485 -205 535 -135
rect 585 -205 635 -190
rect 685 -205 735 -190
rect 785 -205 835 -135
rect 940 -160 980 -150
rect 940 -175 950 -160
rect 885 -180 950 -175
rect 970 -180 980 -160
rect 885 -190 980 -180
rect 885 -205 935 -190
rect -15 -820 35 -805
rect 85 -860 135 -805
rect -95 -870 135 -860
rect 185 -855 235 -805
rect 285 -855 335 -805
rect 385 -820 435 -805
rect 485 -820 535 -805
rect 585 -855 635 -805
rect 685 -855 735 -805
rect 785 -820 835 -805
rect 885 -820 935 -805
rect 185 -865 735 -855
rect 185 -870 450 -865
rect -95 -890 -85 -870
rect -65 -875 135 -870
rect -65 -890 -55 -875
rect -95 -900 -55 -890
rect 440 -885 450 -870
rect 470 -870 735 -865
rect 470 -885 480 -870
rect 440 -895 480 -885
rect 450 -1740 470 -895
rect 380 -1750 540 -1740
rect -60 -1760 -20 -1750
rect -60 -1780 -50 -1760
rect -30 -1775 -20 -1760
rect 380 -1770 390 -1750
rect 410 -1755 510 -1750
rect 410 -1770 420 -1755
rect -30 -1780 100 -1775
rect 380 -1780 420 -1770
rect 500 -1770 510 -1755
rect 530 -1770 540 -1750
rect 500 -1780 540 -1770
rect -60 -1790 100 -1780
rect 85 -1810 100 -1790
rect -60 -1825 -20 -1815
rect -60 -1845 -50 -1825
rect -30 -1840 -20 -1825
rect 85 -1825 835 -1810
rect -30 -1845 35 -1840
rect -60 -1855 35 -1845
rect -15 -1865 35 -1855
rect 85 -1865 135 -1825
rect 185 -1865 235 -1850
rect 285 -1865 335 -1850
rect 385 -1865 435 -1825
rect 485 -1865 535 -1825
rect 585 -1865 635 -1850
rect 685 -1865 735 -1850
rect 785 -1865 835 -1825
rect 940 -1825 980 -1815
rect 940 -1840 950 -1825
rect 885 -1845 950 -1840
rect 970 -1845 980 -1825
rect 885 -1855 980 -1845
rect 885 -1865 935 -1855
rect -15 -2480 35 -2465
rect 85 -2480 135 -2465
rect 185 -2500 235 -2465
rect 285 -2500 335 -2465
rect 385 -2480 435 -2465
rect 485 -2480 535 -2465
rect -65 -2505 -25 -2500
rect 185 -2505 335 -2500
rect 585 -2505 635 -2465
rect 685 -2505 735 -2465
rect 785 -2480 835 -2465
rect 885 -2480 935 -2465
rect -65 -2510 735 -2505
rect -65 -2530 -55 -2510
rect -35 -2520 735 -2510
rect -35 -2530 -25 -2520
rect -65 -2540 -25 -2530
<< polycont >>
rect 95 750 115 770
rect -50 530 -30 550
rect 950 530 970 550
rect 895 455 915 475
rect -50 400 -30 420
rect 950 400 970 420
rect 895 5 915 25
rect 250 -35 270 -15
rect 650 -35 670 -15
rect -50 -180 -30 -160
rect 950 -180 970 -160
rect -85 -890 -65 -870
rect 450 -885 470 -865
rect -50 -1780 -30 -1760
rect 390 -1770 410 -1750
rect 510 -1770 530 -1750
rect -50 -1845 -30 -1825
rect 950 -1845 970 -1825
rect -55 -2530 -35 -2510
<< locali >>
rect 85 770 135 780
rect -115 750 95 770
rect 115 750 135 770
rect 85 745 135 750
rect -110 715 -20 720
rect -110 590 -100 715
rect -80 590 -50 715
rect -30 590 -20 715
rect -110 580 -20 590
rect 40 715 80 720
rect 40 590 50 715
rect 70 590 80 715
rect 40 580 80 590
rect 140 715 180 720
rect 140 590 150 715
rect 170 590 180 715
rect -60 550 -20 580
rect -60 530 -50 550
rect -30 530 -20 550
rect -60 520 -20 530
rect 140 560 180 590
rect 240 715 280 720
rect 240 590 250 715
rect 270 590 280 715
rect 240 580 280 590
rect 340 715 380 720
rect 340 590 350 715
rect 370 590 380 715
rect 340 560 380 590
rect 440 715 480 720
rect 440 590 450 715
rect 470 590 480 715
rect 440 580 480 590
rect 540 715 580 720
rect 540 590 550 715
rect 570 590 580 715
rect 540 560 580 590
rect 640 715 680 720
rect 640 590 650 715
rect 670 590 680 715
rect 640 580 680 590
rect 740 715 780 720
rect 740 590 750 715
rect 770 590 780 715
rect 740 560 780 590
rect 840 715 880 720
rect 840 590 850 715
rect 870 590 880 715
rect 840 580 880 590
rect 940 715 1030 720
rect 940 590 950 715
rect 970 590 1000 715
rect 1020 590 1030 715
rect 940 580 1030 590
rect 140 540 780 560
rect -60 420 -20 430
rect -60 400 -50 420
rect -30 400 -20 420
rect -60 370 -20 400
rect -110 360 -20 370
rect -110 90 -100 360
rect -80 90 -50 360
rect -30 90 -20 360
rect -110 80 -20 90
rect 40 360 80 370
rect 40 90 50 360
rect 70 90 80 360
rect 40 80 80 90
rect 140 360 180 540
rect 140 90 150 360
rect 170 90 180 360
rect 140 80 180 90
rect 240 360 280 370
rect 240 90 250 360
rect 270 90 280 360
rect 60 -45 80 80
rect 240 -15 280 90
rect 340 360 380 540
rect 340 90 350 360
rect 370 90 380 360
rect 340 80 380 90
rect 440 360 480 370
rect 440 90 450 360
rect 470 90 480 360
rect 440 80 480 90
rect 540 360 580 540
rect 540 90 550 360
rect 570 90 580 360
rect 540 80 580 90
rect 640 360 680 370
rect 640 90 650 360
rect 670 90 680 360
rect 240 -35 250 -15
rect 270 -35 280 -15
rect 240 -45 280 -35
rect 60 -55 100 -45
rect 60 -75 70 -55
rect 90 -65 100 -55
rect 450 -65 470 80
rect 640 -15 680 90
rect 740 360 780 540
rect 940 550 980 580
rect 940 530 950 550
rect 970 530 980 550
rect 940 520 980 530
rect 885 475 925 485
rect 885 455 895 475
rect 915 455 1035 475
rect 885 445 925 455
rect 940 420 980 430
rect 940 400 950 420
rect 970 400 980 420
rect 940 370 980 400
rect 740 90 750 360
rect 770 90 780 360
rect 740 80 780 90
rect 840 360 880 370
rect 840 90 850 360
rect 870 90 880 360
rect 840 80 880 90
rect 940 360 1030 370
rect 940 90 950 360
rect 970 90 1000 360
rect 1020 90 1030 360
rect 940 80 1030 90
rect 640 -35 650 -15
rect 670 -35 680 -15
rect 640 -45 680 -35
rect 840 -65 860 80
rect 885 25 1035 35
rect 885 5 895 25
rect 915 15 1035 25
rect 915 5 925 15
rect 885 -5 925 5
rect 90 -75 860 -65
rect 60 -85 860 -75
rect 140 -150 780 -130
rect -60 -160 -20 -150
rect -60 -180 -50 -160
rect -30 -180 -20 -160
rect -60 -210 -20 -180
rect -110 -220 -20 -210
rect -110 -790 -100 -220
rect -80 -790 -50 -220
rect -30 -790 -20 -220
rect -110 -800 -20 -790
rect 40 -220 80 -210
rect 40 -790 50 -220
rect 70 -790 80 -220
rect -115 -870 -55 -860
rect -115 -880 -85 -870
rect -95 -890 -85 -880
rect -65 -890 -55 -870
rect -95 -900 -55 -890
rect 40 -935 80 -790
rect 140 -220 180 -150
rect 340 -190 580 -170
rect 140 -790 150 -220
rect 170 -790 180 -220
rect 140 -800 180 -790
rect 240 -220 280 -210
rect 240 -790 250 -220
rect 270 -790 280 -220
rect 240 -800 280 -790
rect 340 -220 380 -190
rect 340 -790 350 -220
rect 370 -790 380 -220
rect 340 -800 380 -790
rect 440 -220 480 -210
rect 440 -790 450 -220
rect 470 -790 480 -220
rect 440 -865 480 -790
rect 540 -220 580 -190
rect 540 -790 550 -220
rect 570 -790 580 -220
rect 540 -800 580 -790
rect 640 -220 680 -210
rect 640 -790 650 -220
rect 670 -790 680 -220
rect 640 -800 680 -790
rect 740 -220 780 -150
rect 940 -160 980 -150
rect 940 -180 950 -160
rect 970 -180 980 -160
rect 940 -210 980 -180
rect 740 -790 750 -220
rect 770 -790 780 -220
rect 740 -800 780 -790
rect 840 -220 880 -210
rect 840 -790 850 -220
rect 870 -790 880 -220
rect 440 -885 450 -865
rect 470 -885 480 -865
rect 440 -895 480 -885
rect 840 -935 880 -790
rect 940 -220 1030 -210
rect 940 -790 950 -220
rect 970 -790 1000 -220
rect 1020 -790 1030 -220
rect 940 -800 1030 -790
rect -115 -960 -40 -940
rect 40 -955 1035 -935
rect -60 -1750 -40 -960
rect 40 -1750 420 -1740
rect -60 -1760 -20 -1750
rect -60 -1780 -50 -1760
rect -30 -1780 -20 -1760
rect -60 -1790 -20 -1780
rect 40 -1760 390 -1750
rect -60 -1825 -20 -1815
rect -60 -1845 -50 -1825
rect -30 -1845 -20 -1825
rect -60 -1870 -20 -1845
rect -110 -1880 -20 -1870
rect -110 -2450 -100 -1880
rect -80 -2450 -50 -1880
rect -30 -2450 -20 -1880
rect -110 -2460 -20 -2450
rect 40 -1880 80 -1760
rect 380 -1770 390 -1760
rect 410 -1770 420 -1750
rect 380 -1780 420 -1770
rect 40 -2450 50 -1880
rect 70 -2450 80 -1880
rect 40 -2460 80 -2450
rect 140 -1810 180 -1800
rect 140 -1830 150 -1810
rect 170 -1830 180 -1810
rect 140 -1880 180 -1830
rect 140 -2450 150 -1880
rect 170 -2450 180 -1880
rect -115 -2510 -25 -2500
rect -115 -2520 -55 -2510
rect -65 -2530 -55 -2520
rect -35 -2530 -25 -2510
rect -65 -2540 -25 -2530
rect 140 -2520 180 -2450
rect 240 -1880 280 -1870
rect 240 -2450 250 -1880
rect 270 -2450 280 -1880
rect 240 -2460 280 -2450
rect 340 -1880 380 -1870
rect 340 -2450 350 -1880
rect 370 -2450 380 -1880
rect 340 -2480 380 -2450
rect 440 -1880 480 -955
rect 500 -1750 880 -1740
rect 500 -1770 510 -1750
rect 530 -1760 880 -1750
rect 530 -1770 540 -1760
rect 500 -1780 540 -1770
rect 440 -2450 450 -1880
rect 470 -2450 480 -1880
rect 440 -2460 480 -2450
rect 540 -1810 580 -1800
rect 540 -1830 550 -1810
rect 570 -1830 580 -1810
rect 540 -1880 580 -1830
rect 540 -2450 550 -1880
rect 570 -2450 580 -1880
rect 540 -2480 580 -2450
rect 640 -1880 680 -1870
rect 640 -2450 650 -1880
rect 670 -2450 680 -1880
rect 640 -2460 680 -2450
rect 740 -1880 780 -1870
rect 740 -2450 750 -1880
rect 770 -2450 780 -1880
rect 340 -2500 580 -2480
rect 740 -2520 780 -2450
rect 840 -1880 880 -1760
rect 840 -2450 850 -1880
rect 870 -2450 880 -1880
rect 840 -2460 880 -2450
rect 940 -1825 980 -1815
rect 940 -1845 950 -1825
rect 970 -1845 980 -1825
rect 940 -1870 980 -1845
rect 940 -1880 1030 -1870
rect 940 -2450 950 -1880
rect 970 -2450 1000 -1880
rect 1020 -2450 1030 -1880
rect 940 -2460 1030 -2450
rect 140 -2540 780 -2520
<< viali >>
rect -100 590 -80 715
rect -50 590 -30 715
rect 50 590 70 715
rect 250 590 270 715
rect 450 590 470 715
rect 650 590 670 715
rect 850 590 870 715
rect 950 590 970 715
rect 1000 590 1020 715
rect -100 90 -80 360
rect -50 90 -30 360
rect 70 -75 90 -55
rect 950 90 970 360
rect 1000 90 1020 360
rect 650 -35 670 -15
rect -100 -790 -80 -220
rect -50 -790 -30 -220
rect 250 -790 270 -220
rect 650 -790 670 -220
rect 950 -790 970 -220
rect 1000 -790 1020 -220
rect -100 -2450 -80 -1880
rect -50 -2450 -30 -1880
rect 150 -1830 170 -1810
rect 250 -2450 270 -1880
rect 550 -1830 570 -1810
rect 650 -2450 670 -1880
rect 950 -2450 970 -1880
rect 1000 -2450 1020 -1880
<< metal1 >>
rect -115 715 1035 720
rect -115 590 -100 715
rect -80 590 -50 715
rect -30 590 50 715
rect 70 590 250 715
rect 270 590 450 715
rect 470 590 650 715
rect 670 590 850 715
rect 870 590 950 715
rect 970 590 1000 715
rect 1020 590 1035 715
rect -115 360 1035 590
rect -115 90 -100 360
rect -80 90 -50 360
rect -30 90 950 360
rect 970 90 1000 360
rect 1020 90 1035 360
rect -115 80 1035 90
rect -115 -210 -15 80
rect 540 -15 680 -5
rect 540 -35 650 -15
rect 670 -35 680 -15
rect 540 -45 680 -35
rect 60 -55 380 -45
rect 60 -75 70 -55
rect 90 -75 380 -55
rect 60 -85 380 -75
rect -115 -220 280 -210
rect -115 -790 -100 -220
rect -80 -790 -50 -220
rect -30 -790 250 -220
rect 270 -790 280 -220
rect -115 -800 280 -790
rect 340 -1800 380 -85
rect 140 -1810 380 -1800
rect 140 -1830 150 -1810
rect 170 -1830 380 -1810
rect 140 -1840 380 -1830
rect 540 -1810 580 -45
rect 935 -210 1035 80
rect 640 -220 1035 -210
rect 640 -790 650 -220
rect 670 -790 950 -220
rect 970 -790 1000 -220
rect 1020 -790 1035 -220
rect 640 -800 1035 -790
rect 540 -1830 550 -1810
rect 570 -1830 580 -1810
rect 540 -1840 580 -1830
rect -115 -1880 1035 -1870
rect -115 -2450 -100 -1880
rect -80 -2450 -50 -1880
rect -30 -2450 250 -1880
rect 270 -2450 650 -1880
rect 670 -2450 950 -1880
rect 970 -2450 1000 -1880
rect 1020 -2450 1035 -1880
rect -115 -2460 1035 -2450
<< labels >>
rlabel locali -115 -2510 -115 -2510 7 Vbn
rlabel metal1 -115 -2170 -115 -2170 7 Vn
rlabel locali 1035 25 1035 25 3 V2
rlabel locali 1035 465 1035 465 3 V1
rlabel metal1 -115 650 -115 650 7 Vp
rlabel locali -115 760 -115 760 7 Vbp
rlabel locali -115 -870 -115 -870 7 Vcp
rlabel locali -115 -950 -115 -950 7 Vcn
rlabel locali 1035 -945 1035 -945 3 Vout
<< end >>
